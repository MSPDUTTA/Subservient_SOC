VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO subservient
  CLASS BLOCK ;
  FOREIGN subservient ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN i_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 596.000 11.870 600.000 ;
    END
  END i_clk
  PIN i_debug_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END i_debug_mode
  PIN i_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 596.000 34.870 600.000 ;
    END
  END i_rst
  PIN i_sram_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END i_sram_rdata[0]
  PIN i_sram_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END i_sram_rdata[1]
  PIN i_sram_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END i_sram_rdata[2]
  PIN i_sram_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 180.920 900.000 181.520 ;
    END
  END i_sram_rdata[3]
  PIN i_sram_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 227.840 900.000 228.440 ;
    END
  END i_sram_rdata[4]
  PIN i_sram_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.510 596.000 334.790 600.000 ;
    END
  END i_sram_rdata[5]
  PIN i_sram_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END i_sram_rdata[6]
  PIN i_sram_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.000 4.000 202.600 ;
    END
  END i_sram_rdata[7]
  PIN i_wb_dbg_adr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 54.440 900.000 55.040 ;
    END
  END i_wb_dbg_adr[0]
  PIN i_wb_dbg_adr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 323.040 900.000 323.640 ;
    END
  END i_wb_dbg_adr[10]
  PIN i_wb_dbg_adr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 354.320 900.000 354.920 ;
    END
  END i_wb_dbg_adr[11]
  PIN i_wb_dbg_adr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 369.960 900.000 370.560 ;
    END
  END i_wb_dbg_adr[12]
  PIN i_wb_dbg_adr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END i_wb_dbg_adr[13]
  PIN i_wb_dbg_adr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 433.200 900.000 433.800 ;
    END
  END i_wb_dbg_adr[14]
  PIN i_wb_dbg_adr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 465.160 900.000 465.760 ;
    END
  END i_wb_dbg_adr[15]
  PIN i_wb_dbg_adr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END i_wb_dbg_adr[16]
  PIN i_wb_dbg_adr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.280 4.000 369.880 ;
    END
  END i_wb_dbg_adr[17]
  PIN i_wb_dbg_adr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.760 4.000 411.360 ;
    END
  END i_wb_dbg_adr[18]
  PIN i_wb_dbg_adr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END i_wb_dbg_adr[19]
  PIN i_wb_dbg_adr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 596.000 173.330 600.000 ;
    END
  END i_wb_dbg_adr[1]
  PIN i_wb_dbg_adr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 512.080 900.000 512.680 ;
    END
  END i_wb_dbg_adr[20]
  PIN i_wb_dbg_adr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 596.000 634.710 600.000 ;
    END
  END i_wb_dbg_adr[21]
  PIN i_wb_dbg_adr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.470 0.000 645.750 4.000 ;
    END
  END i_wb_dbg_adr[22]
  PIN i_wb_dbg_adr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.890 596.000 727.170 600.000 ;
    END
  END i_wb_dbg_adr[23]
  PIN i_wb_dbg_adr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 596.000 750.170 600.000 ;
    END
  END i_wb_dbg_adr[24]
  PIN i_wb_dbg_adr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 596.000 773.170 600.000 ;
    END
  END i_wb_dbg_adr[25]
  PIN i_wb_dbg_adr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 590.960 900.000 591.560 ;
    END
  END i_wb_dbg_adr[26]
  PIN i_wb_dbg_adr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.770 0.000 763.050 4.000 ;
    END
  END i_wb_dbg_adr[27]
  PIN i_wb_dbg_adr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 522.280 4.000 522.880 ;
    END
  END i_wb_dbg_adr[28]
  PIN i_wb_dbg_adr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.350 596.000 819.630 600.000 ;
    END
  END i_wb_dbg_adr[29]
  PIN i_wb_dbg_adr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 596.000 219.330 600.000 ;
    END
  END i_wb_dbg_adr[2]
  PIN i_wb_dbg_adr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END i_wb_dbg_adr[30]
  PIN i_wb_dbg_adr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.350 596.000 842.630 600.000 ;
    END
  END i_wb_dbg_adr[31]
  PIN i_wb_dbg_adr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END i_wb_dbg_adr[3]
  PIN i_wb_dbg_adr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 596.000 288.790 600.000 ;
    END
  END i_wb_dbg_adr[4]
  PIN i_wb_dbg_adr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END i_wb_dbg_adr[5]
  PIN i_wb_dbg_adr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END i_wb_dbg_adr[6]
  PIN i_wb_dbg_adr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 596.000 450.250 600.000 ;
    END
  END i_wb_dbg_adr[7]
  PIN i_wb_dbg_adr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END i_wb_dbg_adr[8]
  PIN i_wb_dbg_adr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.760 4.000 258.360 ;
    END
  END i_wb_dbg_adr[9]
  PIN i_wb_dbg_dat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 596.000 80.870 600.000 ;
    END
  END i_wb_dbg_dat[0]
  PIN i_wb_dbg_dat[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 338.680 900.000 339.280 ;
    END
  END i_wb_dbg_dat[10]
  PIN i_wb_dbg_dat[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.070 0.000 489.350 4.000 ;
    END
  END i_wb_dbg_dat[11]
  PIN i_wb_dbg_dat[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 313.520 4.000 314.120 ;
    END
  END i_wb_dbg_dat[12]
  PIN i_wb_dbg_dat[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 401.920 900.000 402.520 ;
    END
  END i_wb_dbg_dat[13]
  PIN i_wb_dbg_dat[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 448.840 900.000 449.440 ;
    END
  END i_wb_dbg_dat[14]
  PIN i_wb_dbg_dat[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.430 596.000 588.710 600.000 ;
    END
  END i_wb_dbg_dat[15]
  PIN i_wb_dbg_dat[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END i_wb_dbg_dat[16]
  PIN i_wb_dbg_dat[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.880 4.000 383.480 ;
    END
  END i_wb_dbg_dat[17]
  PIN i_wb_dbg_dat[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END i_wb_dbg_dat[18]
  PIN i_wb_dbg_dat[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END i_wb_dbg_dat[19]
  PIN i_wb_dbg_dat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 596.000 196.330 600.000 ;
    END
  END i_wb_dbg_dat[1]
  PIN i_wb_dbg_dat[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 527.720 900.000 528.320 ;
    END
  END i_wb_dbg_dat[20]
  PIN i_wb_dbg_dat[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.890 596.000 658.170 600.000 ;
    END
  END i_wb_dbg_dat[21]
  PIN i_wb_dbg_dat[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.890 596.000 681.170 600.000 ;
    END
  END i_wb_dbg_dat[22]
  PIN i_wb_dbg_dat[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 559.680 900.000 560.280 ;
    END
  END i_wb_dbg_dat[23]
  PIN i_wb_dbg_dat[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.800 4.000 481.400 ;
    END
  END i_wb_dbg_dat[24]
  PIN i_wb_dbg_dat[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 494.400 4.000 495.000 ;
    END
  END i_wb_dbg_dat[25]
  PIN i_wb_dbg_dat[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.670 0.000 723.950 4.000 ;
    END
  END i_wb_dbg_dat[26]
  PIN i_wb_dbg_dat[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.350 596.000 796.630 600.000 ;
    END
  END i_wb_dbg_dat[27]
  PIN i_wb_dbg_dat[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 536.560 4.000 537.160 ;
    END
  END i_wb_dbg_dat[28]
  PIN i_wb_dbg_dat[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END i_wb_dbg_dat[29]
  PIN i_wb_dbg_dat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END i_wb_dbg_dat[2]
  PIN i_wb_dbg_dat[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.070 0.000 880.350 4.000 ;
    END
  END i_wb_dbg_dat[30]
  PIN i_wb_dbg_dat[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.350 596.000 865.630 600.000 ;
    END
  END i_wb_dbg_dat[31]
  PIN i_wb_dbg_dat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 196.560 900.000 197.160 ;
    END
  END i_wb_dbg_dat[3]
  PIN i_wb_dbg_dat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 596.000 311.790 600.000 ;
    END
  END i_wb_dbg_dat[4]
  PIN i_wb_dbg_dat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 275.440 900.000 276.040 ;
    END
  END i_wb_dbg_dat[5]
  PIN i_wb_dbg_dat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 596.000 404.250 600.000 ;
    END
  END i_wb_dbg_dat[6]
  PIN i_wb_dbg_dat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 291.080 900.000 291.680 ;
    END
  END i_wb_dbg_dat[7]
  PIN i_wb_dbg_dat[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 307.400 900.000 308.000 ;
    END
  END i_wb_dbg_dat[8]
  PIN i_wb_dbg_dat[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.430 596.000 565.710 600.000 ;
    END
  END i_wb_dbg_dat[9]
  PIN i_wb_dbg_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 596.000 103.870 600.000 ;
    END
  END i_wb_dbg_sel[0]
  PIN i_wb_dbg_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 102.040 900.000 102.640 ;
    END
  END i_wb_dbg_sel[1]
  PIN i_wb_dbg_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 148.960 900.000 149.560 ;
    END
  END i_wb_dbg_sel[2]
  PIN i_wb_dbg_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 0.000 215.190 4.000 ;
    END
  END i_wb_dbg_sel[3]
  PIN i_wb_dbg_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 7.520 900.000 8.120 ;
    END
  END i_wb_dbg_stb
  PIN i_wb_dbg_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 596.000 57.870 600.000 ;
    END
  END i_wb_dbg_we
  PIN o_gpio
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 23.160 900.000 23.760 ;
    END
  END o_gpio
  PIN o_sram_raddr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 70.080 900.000 70.680 ;
    END
  END o_sram_raddr[0]
  PIN o_sram_raddr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 117.680 900.000 118.280 ;
    END
  END o_sram_raddr[1]
  PIN o_sram_raddr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 165.280 900.000 165.880 ;
    END
  END o_sram_raddr[2]
  PIN o_sram_raddr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 596.000 242.330 600.000 ;
    END
  END o_sram_raddr[3]
  PIN o_sram_raddr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END o_sram_raddr[4]
  PIN o_sram_raddr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END o_sram_raddr[5]
  PIN o_sram_raddr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 0.000 371.590 4.000 ;
    END
  END o_sram_raddr[6]
  PIN o_sram_raddr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.600 4.000 216.200 ;
    END
  END o_sram_raddr[7]
  PIN o_sram_raddr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.970 596.000 519.250 600.000 ;
    END
  END o_sram_raddr[8]
  PIN o_sram_ren
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END o_sram_ren
  PIN o_sram_waddr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 86.400 900.000 87.000 ;
    END
  END o_sram_waddr[0]
  PIN o_sram_waddr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 133.320 900.000 133.920 ;
    END
  END o_sram_waddr[1]
  PIN o_sram_waddr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END o_sram_waddr[2]
  PIN o_sram_waddr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 212.200 900.000 212.800 ;
    END
  END o_sram_waddr[3]
  PIN o_sram_waddr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 244.160 900.000 244.760 ;
    END
  END o_sram_waddr[4]
  PIN o_sram_waddr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 596.000 357.790 600.000 ;
    END
  END o_sram_waddr[5]
  PIN o_sram_waddr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.970 596.000 427.250 600.000 ;
    END
  END o_sram_waddr[6]
  PIN o_sram_waddr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END o_sram_waddr[7]
  PIN o_sram_waddr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END o_sram_waddr[8]
  PIN o_sram_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 596.000 126.870 600.000 ;
    END
  END o_sram_wdata[0]
  PIN o_sram_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END o_sram_wdata[1]
  PIN o_sram_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END o_sram_wdata[2]
  PIN o_sram_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 596.000 265.330 600.000 ;
    END
  END o_sram_wdata[3]
  PIN o_sram_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 259.800 900.000 260.400 ;
    END
  END o_sram_wdata[4]
  PIN o_sram_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END o_sram_wdata[5]
  PIN o_sram_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END o_sram_wdata[6]
  PIN o_sram_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.970 596.000 473.250 600.000 ;
    END
  END o_sram_wdata[7]
  PIN o_sram_wen
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 38.800 900.000 39.400 ;
    END
  END o_sram_wen
  PIN o_wb_dbg_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END o_wb_dbg_ack
  PIN o_wb_dbg_rdt[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 596.000 150.330 600.000 ;
    END
  END o_wb_dbg_rdt[0]
  PIN o_wb_dbg_rdt[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END o_wb_dbg_rdt[10]
  PIN o_wb_dbg_rdt[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END o_wb_dbg_rdt[11]
  PIN o_wb_dbg_rdt[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 386.280 900.000 386.880 ;
    END
  END o_wb_dbg_rdt[12]
  PIN o_wb_dbg_rdt[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 417.560 900.000 418.160 ;
    END
  END o_wb_dbg_rdt[13]
  PIN o_wb_dbg_rdt[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 0.000 567.550 4.000 ;
    END
  END o_wb_dbg_rdt[14]
  PIN o_wb_dbg_rdt[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.120 4.000 327.720 ;
    END
  END o_wb_dbg_rdt[15]
  PIN o_wb_dbg_rdt[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 480.800 900.000 481.400 ;
    END
  END o_wb_dbg_rdt[16]
  PIN o_wb_dbg_rdt[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END o_wb_dbg_rdt[17]
  PIN o_wb_dbg_rdt[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 496.440 900.000 497.040 ;
    END
  END o_wb_dbg_rdt[18]
  PIN o_wb_dbg_rdt[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.370 0.000 606.650 4.000 ;
    END
  END o_wb_dbg_rdt[19]
  PIN o_wb_dbg_rdt[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 4.000 91.080 ;
    END
  END o_wb_dbg_rdt[1]
  PIN o_wb_dbg_rdt[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.430 596.000 611.710 600.000 ;
    END
  END o_wb_dbg_rdt[20]
  PIN o_wb_dbg_rdt[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 544.040 900.000 544.640 ;
    END
  END o_wb_dbg_rdt[21]
  PIN o_wb_dbg_rdt[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 596.000 704.170 600.000 ;
    END
  END o_wb_dbg_rdt[22]
  PIN o_wb_dbg_rdt[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.520 4.000 467.120 ;
    END
  END o_wb_dbg_rdt[23]
  PIN o_wb_dbg_rdt[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.570 0.000 684.850 4.000 ;
    END
  END o_wb_dbg_rdt[24]
  PIN o_wb_dbg_rdt[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 575.320 900.000 575.920 ;
    END
  END o_wb_dbg_rdt[25]
  PIN o_wb_dbg_rdt[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.680 4.000 509.280 ;
    END
  END o_wb_dbg_rdt[26]
  PIN o_wb_dbg_rdt[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 0.000 802.150 4.000 ;
    END
  END o_wb_dbg_rdt[27]
  PIN o_wb_dbg_rdt[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.160 4.000 550.760 ;
    END
  END o_wb_dbg_rdt[28]
  PIN o_wb_dbg_rdt[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.970 0.000 841.250 4.000 ;
    END
  END o_wb_dbg_rdt[29]
  PIN o_wb_dbg_rdt[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.080 4.000 104.680 ;
    END
  END o_wb_dbg_rdt[2]
  PIN o_wb_dbg_rdt[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 592.320 4.000 592.920 ;
    END
  END o_wb_dbg_rdt[30]
  PIN o_wb_dbg_rdt[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.350 596.000 888.630 600.000 ;
    END
  END o_wb_dbg_rdt[31]
  PIN o_wb_dbg_rdt[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END o_wb_dbg_rdt[3]
  PIN o_wb_dbg_rdt[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END o_wb_dbg_rdt[4]
  PIN o_wb_dbg_rdt[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 596.000 380.790 600.000 ;
    END
  END o_wb_dbg_rdt[5]
  PIN o_wb_dbg_rdt[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 0.000 410.690 4.000 ;
    END
  END o_wb_dbg_rdt[6]
  PIN o_wb_dbg_rdt[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 596.000 496.250 600.000 ;
    END
  END o_wb_dbg_rdt[7]
  PIN o_wb_dbg_rdt[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 596.000 542.710 600.000 ;
    END
  END o_wb_dbg_rdt[8]
  PIN o_wb_dbg_rdt[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 271.360 4.000 271.960 ;
    END
  END o_wb_dbg_rdt[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 792.340 10.880 793.940 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 638.740 10.880 640.340 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 485.140 10.880 486.740 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.540 10.880 333.140 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 587.520 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 869.140 10.880 870.740 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 715.540 10.880 717.140 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 561.940 10.880 563.540 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 408.340 10.880 409.940 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.740 10.880 256.340 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 587.520 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 795.640 10.880 797.240 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 642.040 10.880 643.640 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 488.440 10.880 490.040 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 334.840 10.880 336.440 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.240 10.880 182.840 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.640 10.880 29.240 587.520 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 872.440 10.880 874.040 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 718.840 10.880 720.440 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 565.240 10.880 566.840 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 411.640 10.880 413.240 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 258.040 10.880 259.640 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.440 10.880 106.040 587.520 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 798.940 10.880 800.540 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 645.340 10.880 646.940 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 491.740 10.880 493.340 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 338.140 10.880 339.740 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.540 10.880 186.140 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.880 32.540 587.520 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 875.740 10.880 877.340 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 722.140 10.880 723.740 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 568.540 10.880 570.140 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 414.940 10.880 416.540 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 261.340 10.880 262.940 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.740 10.880 109.340 587.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 894.240 587.605 ;
      LAYER met1 ;
        RECT 5.520 10.640 894.240 587.760 ;
      LAYER met2 ;
        RECT 10.210 595.720 11.310 596.000 ;
        RECT 12.150 595.720 34.310 596.000 ;
        RECT 35.150 595.720 57.310 596.000 ;
        RECT 58.150 595.720 80.310 596.000 ;
        RECT 81.150 595.720 103.310 596.000 ;
        RECT 104.150 595.720 126.310 596.000 ;
        RECT 127.150 595.720 149.770 596.000 ;
        RECT 150.610 595.720 172.770 596.000 ;
        RECT 173.610 595.720 195.770 596.000 ;
        RECT 196.610 595.720 218.770 596.000 ;
        RECT 219.610 595.720 241.770 596.000 ;
        RECT 242.610 595.720 264.770 596.000 ;
        RECT 265.610 595.720 288.230 596.000 ;
        RECT 289.070 595.720 311.230 596.000 ;
        RECT 312.070 595.720 334.230 596.000 ;
        RECT 335.070 595.720 357.230 596.000 ;
        RECT 358.070 595.720 380.230 596.000 ;
        RECT 381.070 595.720 403.690 596.000 ;
        RECT 404.530 595.720 426.690 596.000 ;
        RECT 427.530 595.720 449.690 596.000 ;
        RECT 450.530 595.720 472.690 596.000 ;
        RECT 473.530 595.720 495.690 596.000 ;
        RECT 496.530 595.720 518.690 596.000 ;
        RECT 519.530 595.720 542.150 596.000 ;
        RECT 542.990 595.720 565.150 596.000 ;
        RECT 565.990 595.720 588.150 596.000 ;
        RECT 588.990 595.720 611.150 596.000 ;
        RECT 611.990 595.720 634.150 596.000 ;
        RECT 634.990 595.720 657.610 596.000 ;
        RECT 658.450 595.720 680.610 596.000 ;
        RECT 681.450 595.720 703.610 596.000 ;
        RECT 704.450 595.720 726.610 596.000 ;
        RECT 727.450 595.720 749.610 596.000 ;
        RECT 750.450 595.720 772.610 596.000 ;
        RECT 773.450 595.720 796.070 596.000 ;
        RECT 796.910 595.720 819.070 596.000 ;
        RECT 819.910 595.720 842.070 596.000 ;
        RECT 842.910 595.720 865.070 596.000 ;
        RECT 865.910 595.720 888.070 596.000 ;
        RECT 10.210 4.280 888.620 595.720 ;
        RECT 10.210 4.000 19.130 4.280 ;
        RECT 19.970 4.000 58.230 4.280 ;
        RECT 59.070 4.000 97.330 4.280 ;
        RECT 98.170 4.000 136.430 4.280 ;
        RECT 137.270 4.000 175.530 4.280 ;
        RECT 176.370 4.000 214.630 4.280 ;
        RECT 215.470 4.000 253.730 4.280 ;
        RECT 254.570 4.000 292.830 4.280 ;
        RECT 293.670 4.000 331.930 4.280 ;
        RECT 332.770 4.000 371.030 4.280 ;
        RECT 371.870 4.000 410.130 4.280 ;
        RECT 410.970 4.000 449.230 4.280 ;
        RECT 450.070 4.000 488.790 4.280 ;
        RECT 489.630 4.000 527.890 4.280 ;
        RECT 528.730 4.000 566.990 4.280 ;
        RECT 567.830 4.000 606.090 4.280 ;
        RECT 606.930 4.000 645.190 4.280 ;
        RECT 646.030 4.000 684.290 4.280 ;
        RECT 685.130 4.000 723.390 4.280 ;
        RECT 724.230 4.000 762.490 4.280 ;
        RECT 763.330 4.000 801.590 4.280 ;
        RECT 802.430 4.000 840.690 4.280 ;
        RECT 841.530 4.000 879.790 4.280 ;
        RECT 880.630 4.000 888.620 4.280 ;
      LAYER met3 ;
        RECT 4.400 591.960 896.000 592.785 ;
        RECT 4.400 591.920 895.600 591.960 ;
        RECT 4.000 590.560 895.600 591.920 ;
        RECT 4.000 579.040 896.000 590.560 ;
        RECT 4.400 577.640 896.000 579.040 ;
        RECT 4.000 576.320 896.000 577.640 ;
        RECT 4.000 574.920 895.600 576.320 ;
        RECT 4.000 565.440 896.000 574.920 ;
        RECT 4.400 564.040 896.000 565.440 ;
        RECT 4.000 560.680 896.000 564.040 ;
        RECT 4.000 559.280 895.600 560.680 ;
        RECT 4.000 551.160 896.000 559.280 ;
        RECT 4.400 549.760 896.000 551.160 ;
        RECT 4.000 545.040 896.000 549.760 ;
        RECT 4.000 543.640 895.600 545.040 ;
        RECT 4.000 537.560 896.000 543.640 ;
        RECT 4.400 536.160 896.000 537.560 ;
        RECT 4.000 528.720 896.000 536.160 ;
        RECT 4.000 527.320 895.600 528.720 ;
        RECT 4.000 523.280 896.000 527.320 ;
        RECT 4.400 521.880 896.000 523.280 ;
        RECT 4.000 513.080 896.000 521.880 ;
        RECT 4.000 511.680 895.600 513.080 ;
        RECT 4.000 509.680 896.000 511.680 ;
        RECT 4.400 508.280 896.000 509.680 ;
        RECT 4.000 497.440 896.000 508.280 ;
        RECT 4.000 496.040 895.600 497.440 ;
        RECT 4.000 495.400 896.000 496.040 ;
        RECT 4.400 494.000 896.000 495.400 ;
        RECT 4.000 481.800 896.000 494.000 ;
        RECT 4.400 480.400 895.600 481.800 ;
        RECT 4.000 467.520 896.000 480.400 ;
        RECT 4.400 466.160 896.000 467.520 ;
        RECT 4.400 466.120 895.600 466.160 ;
        RECT 4.000 464.760 895.600 466.120 ;
        RECT 4.000 453.920 896.000 464.760 ;
        RECT 4.400 452.520 896.000 453.920 ;
        RECT 4.000 449.840 896.000 452.520 ;
        RECT 4.000 448.440 895.600 449.840 ;
        RECT 4.000 439.640 896.000 448.440 ;
        RECT 4.400 438.240 896.000 439.640 ;
        RECT 4.000 434.200 896.000 438.240 ;
        RECT 4.000 432.800 895.600 434.200 ;
        RECT 4.000 426.040 896.000 432.800 ;
        RECT 4.400 424.640 896.000 426.040 ;
        RECT 4.000 418.560 896.000 424.640 ;
        RECT 4.000 417.160 895.600 418.560 ;
        RECT 4.000 411.760 896.000 417.160 ;
        RECT 4.400 410.360 896.000 411.760 ;
        RECT 4.000 402.920 896.000 410.360 ;
        RECT 4.000 401.520 895.600 402.920 ;
        RECT 4.000 398.160 896.000 401.520 ;
        RECT 4.400 396.760 896.000 398.160 ;
        RECT 4.000 387.280 896.000 396.760 ;
        RECT 4.000 385.880 895.600 387.280 ;
        RECT 4.000 383.880 896.000 385.880 ;
        RECT 4.400 382.480 896.000 383.880 ;
        RECT 4.000 370.960 896.000 382.480 ;
        RECT 4.000 370.280 895.600 370.960 ;
        RECT 4.400 369.560 895.600 370.280 ;
        RECT 4.400 368.880 896.000 369.560 ;
        RECT 4.000 356.000 896.000 368.880 ;
        RECT 4.400 355.320 896.000 356.000 ;
        RECT 4.400 354.600 895.600 355.320 ;
        RECT 4.000 353.920 895.600 354.600 ;
        RECT 4.000 342.400 896.000 353.920 ;
        RECT 4.400 341.000 896.000 342.400 ;
        RECT 4.000 339.680 896.000 341.000 ;
        RECT 4.000 338.280 895.600 339.680 ;
        RECT 4.000 328.120 896.000 338.280 ;
        RECT 4.400 326.720 896.000 328.120 ;
        RECT 4.000 324.040 896.000 326.720 ;
        RECT 4.000 322.640 895.600 324.040 ;
        RECT 4.000 314.520 896.000 322.640 ;
        RECT 4.400 313.120 896.000 314.520 ;
        RECT 4.000 308.400 896.000 313.120 ;
        RECT 4.000 307.000 895.600 308.400 ;
        RECT 4.000 300.240 896.000 307.000 ;
        RECT 4.400 298.840 896.000 300.240 ;
        RECT 4.000 292.080 896.000 298.840 ;
        RECT 4.000 290.680 895.600 292.080 ;
        RECT 4.000 286.640 896.000 290.680 ;
        RECT 4.400 285.240 896.000 286.640 ;
        RECT 4.000 276.440 896.000 285.240 ;
        RECT 4.000 275.040 895.600 276.440 ;
        RECT 4.000 272.360 896.000 275.040 ;
        RECT 4.400 270.960 896.000 272.360 ;
        RECT 4.000 260.800 896.000 270.960 ;
        RECT 4.000 259.400 895.600 260.800 ;
        RECT 4.000 258.760 896.000 259.400 ;
        RECT 4.400 257.360 896.000 258.760 ;
        RECT 4.000 245.160 896.000 257.360 ;
        RECT 4.000 244.480 895.600 245.160 ;
        RECT 4.400 243.760 895.600 244.480 ;
        RECT 4.400 243.080 896.000 243.760 ;
        RECT 4.000 230.880 896.000 243.080 ;
        RECT 4.400 229.480 896.000 230.880 ;
        RECT 4.000 228.840 896.000 229.480 ;
        RECT 4.000 227.440 895.600 228.840 ;
        RECT 4.000 216.600 896.000 227.440 ;
        RECT 4.400 215.200 896.000 216.600 ;
        RECT 4.000 213.200 896.000 215.200 ;
        RECT 4.000 211.800 895.600 213.200 ;
        RECT 4.000 203.000 896.000 211.800 ;
        RECT 4.400 201.600 896.000 203.000 ;
        RECT 4.000 197.560 896.000 201.600 ;
        RECT 4.000 196.160 895.600 197.560 ;
        RECT 4.000 188.720 896.000 196.160 ;
        RECT 4.400 187.320 896.000 188.720 ;
        RECT 4.000 181.920 896.000 187.320 ;
        RECT 4.000 180.520 895.600 181.920 ;
        RECT 4.000 175.120 896.000 180.520 ;
        RECT 4.400 173.720 896.000 175.120 ;
        RECT 4.000 166.280 896.000 173.720 ;
        RECT 4.000 164.880 895.600 166.280 ;
        RECT 4.000 160.840 896.000 164.880 ;
        RECT 4.400 159.440 896.000 160.840 ;
        RECT 4.000 149.960 896.000 159.440 ;
        RECT 4.000 148.560 895.600 149.960 ;
        RECT 4.000 147.240 896.000 148.560 ;
        RECT 4.400 145.840 896.000 147.240 ;
        RECT 4.000 134.320 896.000 145.840 ;
        RECT 4.000 132.960 895.600 134.320 ;
        RECT 4.400 132.920 895.600 132.960 ;
        RECT 4.400 131.560 896.000 132.920 ;
        RECT 4.000 119.360 896.000 131.560 ;
        RECT 4.400 118.680 896.000 119.360 ;
        RECT 4.400 117.960 895.600 118.680 ;
        RECT 4.000 117.280 895.600 117.960 ;
        RECT 4.000 105.080 896.000 117.280 ;
        RECT 4.400 103.680 896.000 105.080 ;
        RECT 4.000 103.040 896.000 103.680 ;
        RECT 4.000 101.640 895.600 103.040 ;
        RECT 4.000 91.480 896.000 101.640 ;
        RECT 4.400 90.080 896.000 91.480 ;
        RECT 4.000 87.400 896.000 90.080 ;
        RECT 4.000 86.000 895.600 87.400 ;
        RECT 4.000 77.200 896.000 86.000 ;
        RECT 4.400 75.800 896.000 77.200 ;
        RECT 4.000 71.080 896.000 75.800 ;
        RECT 4.000 69.680 895.600 71.080 ;
        RECT 4.000 63.600 896.000 69.680 ;
        RECT 4.400 62.200 896.000 63.600 ;
        RECT 4.000 55.440 896.000 62.200 ;
        RECT 4.000 54.040 895.600 55.440 ;
        RECT 4.000 49.320 896.000 54.040 ;
        RECT 4.400 47.920 896.000 49.320 ;
        RECT 4.000 39.800 896.000 47.920 ;
        RECT 4.000 38.400 895.600 39.800 ;
        RECT 4.000 35.720 896.000 38.400 ;
        RECT 4.400 34.320 896.000 35.720 ;
        RECT 4.000 24.160 896.000 34.320 ;
        RECT 4.000 22.760 895.600 24.160 ;
        RECT 4.000 21.440 896.000 22.760 ;
        RECT 4.400 20.040 896.000 21.440 ;
        RECT 4.000 8.520 896.000 20.040 ;
        RECT 4.000 7.840 895.600 8.520 ;
        RECT 4.400 7.120 895.600 7.840 ;
        RECT 4.400 6.975 896.000 7.120 ;
      LAYER met4 ;
        RECT 340.695 20.575 401.745 311.265 ;
  END
END subservient
END LIBRARY

