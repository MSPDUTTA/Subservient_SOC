VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO subservient
  CLASS BLOCK ;
  FOREIGN subservient ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN i_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 596.000 14.630 600.000 ;
    END
  END i_clk
  PIN i_debug_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 8.200 900.000 8.800 ;
    END
  END i_debug_mode
  PIN i_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END i_rst
  PIN i_sram_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 596.000 130.550 600.000 ;
    END
  END i_sram_rdata[0]
  PIN i_sram_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END i_sram_rdata[1]
  PIN i_sram_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 596.000 246.930 600.000 ;
    END
  END i_sram_rdata[2]
  PIN i_sram_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 124.480 900.000 125.080 ;
    END
  END i_sram_rdata[3]
  PIN i_sram_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 596.000 333.870 600.000 ;
    END
  END i_sram_rdata[4]
  PIN i_sram_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 4.000 ;
    END
  END i_sram_rdata[5]
  PIN i_sram_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END i_sram_rdata[6]
  PIN i_sram_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END i_sram_rdata[7]
  PIN i_wb_dbg_adr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 41.520 900.000 42.120 ;
    END
  END i_wb_dbg_adr[0]
  PIN i_wb_dbg_adr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END i_wb_dbg_adr[10]
  PIN i_wb_dbg_adr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 0.000 427.710 4.000 ;
    END
  END i_wb_dbg_adr[11]
  PIN i_wb_dbg_adr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 324.400 900.000 325.000 ;
    END
  END i_wb_dbg_adr[12]
  PIN i_wb_dbg_adr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.870 596.000 595.150 600.000 ;
    END
  END i_wb_dbg_adr[13]
  PIN i_wb_dbg_adr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 0.000 515.570 4.000 ;
    END
  END i_wb_dbg_adr[14]
  PIN i_wb_dbg_adr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 357.720 900.000 358.320 ;
    END
  END i_wb_dbg_adr[15]
  PIN i_wb_dbg_adr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 453.600 4.000 454.200 ;
    END
  END i_wb_dbg_adr[16]
  PIN i_wb_dbg_adr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.530 0.000 581.810 4.000 ;
    END
  END i_wb_dbg_adr[17]
  PIN i_wb_dbg_adr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.830 596.000 653.110 600.000 ;
    END
  END i_wb_dbg_adr[18]
  PIN i_wb_dbg_adr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 408.040 900.000 408.640 ;
    END
  END i_wb_dbg_adr[19]
  PIN i_wb_dbg_adr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END i_wb_dbg_adr[1]
  PIN i_wb_dbg_adr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 504.600 4.000 505.200 ;
    END
  END i_wb_dbg_adr[20]
  PIN i_wb_dbg_adr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.810 596.000 682.090 600.000 ;
    END
  END i_wb_dbg_adr[21]
  PIN i_wb_dbg_adr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 522.280 4.000 522.880 ;
    END
  END i_wb_dbg_adr[22]
  PIN i_wb_dbg_adr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.250 596.000 711.530 600.000 ;
    END
  END i_wb_dbg_adr[23]
  PIN i_wb_dbg_adr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 441.360 900.000 441.960 ;
    END
  END i_wb_dbg_adr[24]
  PIN i_wb_dbg_adr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.950 0.000 801.230 4.000 ;
    END
  END i_wb_dbg_adr[25]
  PIN i_wb_dbg_adr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 491.000 900.000 491.600 ;
    END
  END i_wb_dbg_adr[26]
  PIN i_wb_dbg_adr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.210 596.000 769.490 600.000 ;
    END
  END i_wb_dbg_adr[27]
  PIN i_wb_dbg_adr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 524.320 900.000 524.920 ;
    END
  END i_wb_dbg_adr[28]
  PIN i_wb_dbg_adr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.730 0.000 867.010 4.000 ;
    END
  END i_wb_dbg_adr[29]
  PIN i_wb_dbg_adr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 108.160 900.000 108.760 ;
    END
  END i_wb_dbg_adr[2]
  PIN i_wb_dbg_adr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 0.000 889.090 4.000 ;
    END
  END i_wb_dbg_adr[30]
  PIN i_wb_dbg_adr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.130 596.000 885.410 600.000 ;
    END
  END i_wb_dbg_adr[31]
  PIN i_wb_dbg_adr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END i_wb_dbg_adr[3]
  PIN i_wb_dbg_adr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 596.000 362.850 600.000 ;
    END
  END i_wb_dbg_adr[4]
  PIN i_wb_dbg_adr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END i_wb_dbg_adr[5]
  PIN i_wb_dbg_adr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 274.760 900.000 275.360 ;
    END
  END i_wb_dbg_adr[6]
  PIN i_wb_dbg_adr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 596.000 449.790 600.000 ;
    END
  END i_wb_dbg_adr[7]
  PIN i_wb_dbg_adr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 291.080 900.000 291.680 ;
    END
  END i_wb_dbg_adr[8]
  PIN i_wb_dbg_adr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END i_wb_dbg_adr[9]
  PIN i_wb_dbg_dat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 596.000 159.530 600.000 ;
    END
  END i_wb_dbg_dat[0]
  PIN i_wb_dbg_dat[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END i_wb_dbg_dat[10]
  PIN i_wb_dbg_dat[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END i_wb_dbg_dat[11]
  PIN i_wb_dbg_dat[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END i_wb_dbg_dat[12]
  PIN i_wb_dbg_dat[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.670 0.000 493.950 4.000 ;
    END
  END i_wb_dbg_dat[13]
  PIN i_wb_dbg_dat[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 341.400 900.000 342.000 ;
    END
  END i_wb_dbg_dat[14]
  PIN i_wb_dbg_dat[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END i_wb_dbg_dat[15]
  PIN i_wb_dbg_dat[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 596.000 624.130 600.000 ;
    END
  END i_wb_dbg_dat[16]
  PIN i_wb_dbg_dat[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 391.040 900.000 391.640 ;
    END
  END i_wb_dbg_dat[17]
  PIN i_wb_dbg_dat[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 487.600 4.000 488.200 ;
    END
  END i_wb_dbg_dat[18]
  PIN i_wb_dbg_dat[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.230 0.000 625.510 4.000 ;
    END
  END i_wb_dbg_dat[19]
  PIN i_wb_dbg_dat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 4.000 111.480 ;
    END
  END i_wb_dbg_dat[1]
  PIN i_wb_dbg_dat[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.930 0.000 669.210 4.000 ;
    END
  END i_wb_dbg_dat[20]
  PIN i_wb_dbg_dat[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.010 0.000 691.290 4.000 ;
    END
  END i_wb_dbg_dat[21]
  PIN i_wb_dbg_dat[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.170 0.000 735.450 4.000 ;
    END
  END i_wb_dbg_dat[22]
  PIN i_wb_dbg_dat[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.870 0.000 779.150 4.000 ;
    END
  END i_wb_dbg_dat[23]
  PIN i_wb_dbg_dat[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.230 596.000 740.510 600.000 ;
    END
  END i_wb_dbg_dat[24]
  PIN i_wb_dbg_dat[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 474.680 900.000 475.280 ;
    END
  END i_wb_dbg_dat[25]
  PIN i_wb_dbg_dat[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.030 0.000 823.310 4.000 ;
    END
  END i_wb_dbg_dat[26]
  PIN i_wb_dbg_dat[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.650 0.000 844.930 4.000 ;
    END
  END i_wb_dbg_dat[27]
  PIN i_wb_dbg_dat[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.190 596.000 798.470 600.000 ;
    END
  END i_wb_dbg_dat[28]
  PIN i_wb_dbg_dat[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.170 596.000 827.450 600.000 ;
    END
  END i_wb_dbg_dat[29]
  PIN i_wb_dbg_dat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END i_wb_dbg_dat[2]
  PIN i_wb_dbg_dat[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 557.640 900.000 558.240 ;
    END
  END i_wb_dbg_dat[30]
  PIN i_wb_dbg_dat[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.280 4.000 590.880 ;
    END
  END i_wb_dbg_dat[31]
  PIN i_wb_dbg_dat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 4.000 ;
    END
  END i_wb_dbg_dat[3]
  PIN i_wb_dbg_dat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 596.000 391.830 600.000 ;
    END
  END i_wb_dbg_dat[4]
  PIN i_wb_dbg_dat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 224.440 900.000 225.040 ;
    END
  END i_wb_dbg_dat[5]
  PIN i_wb_dbg_dat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 4.000 ;
    END
  END i_wb_dbg_dat[6]
  PIN i_wb_dbg_dat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 596.000 479.230 600.000 ;
    END
  END i_wb_dbg_dat[7]
  PIN i_wb_dbg_dat[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END i_wb_dbg_dat[8]
  PIN i_wb_dbg_dat[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.890 596.000 566.170 600.000 ;
    END
  END i_wb_dbg_dat[9]
  PIN i_wb_dbg_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 596.000 188.510 600.000 ;
    END
  END i_wb_dbg_sel[0]
  PIN i_wb_dbg_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END i_wb_dbg_sel[1]
  PIN i_wb_dbg_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.880 4.000 145.480 ;
    END
  END i_wb_dbg_sel[2]
  PIN i_wb_dbg_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END i_wb_dbg_sel[3]
  PIN i_wb_dbg_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END i_wb_dbg_stb
  PIN i_wb_dbg_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 596.000 43.610 600.000 ;
    END
  END i_wb_dbg_we
  PIN o_gpio
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 596.000 72.590 600.000 ;
    END
  END o_gpio
  PIN o_sram_raddr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 596.000 217.490 600.000 ;
    END
  END o_sram_raddr[0]
  PIN o_sram_raddr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END o_sram_raddr[1]
  PIN o_sram_raddr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END o_sram_raddr[2]
  PIN o_sram_raddr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 141.480 900.000 142.080 ;
    END
  END o_sram_raddr[3]
  PIN o_sram_raddr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END o_sram_raddr[4]
  PIN o_sram_raddr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 241.440 900.000 242.040 ;
    END
  END o_sram_raddr[5]
  PIN o_sram_raddr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END o_sram_raddr[6]
  PIN o_sram_raddr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.930 596.000 508.210 600.000 ;
    END
  END o_sram_raddr[7]
  PIN o_sram_raddr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 308.080 900.000 308.680 ;
    END
  END o_sram_raddr[8]
  PIN o_sram_ren
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 24.520 900.000 25.120 ;
    END
  END o_sram_ren
  PIN o_sram_waddr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 4.000 ;
    END
  END o_sram_waddr[0]
  PIN o_sram_waddr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END o_sram_waddr[1]
  PIN o_sram_waddr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 596.000 275.910 600.000 ;
    END
  END o_sram_waddr[2]
  PIN o_sram_waddr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END o_sram_waddr[3]
  PIN o_sram_waddr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 191.120 900.000 191.720 ;
    END
  END o_sram_waddr[4]
  PIN o_sram_waddr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END o_sram_waddr[5]
  PIN o_sram_waddr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 4.000 ;
    END
  END o_sram_waddr[6]
  PIN o_sram_waddr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 4.000 ;
    END
  END o_sram_waddr[7]
  PIN o_sram_waddr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.730 0.000 384.010 4.000 ;
    END
  END o_sram_waddr[8]
  PIN o_sram_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END o_sram_wdata[0]
  PIN o_sram_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 74.840 900.000 75.440 ;
    END
  END o_sram_wdata[1]
  PIN o_sram_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END o_sram_wdata[2]
  PIN o_sram_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 157.800 900.000 158.400 ;
    END
  END o_sram_wdata[3]
  PIN o_sram_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 208.120 900.000 208.720 ;
    END
  END o_sram_wdata[4]
  PIN o_sram_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 257.760 900.000 258.360 ;
    END
  END o_sram_wdata[5]
  PIN o_sram_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 230.560 4.000 231.160 ;
    END
  END o_sram_wdata[6]
  PIN o_sram_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END o_sram_wdata[7]
  PIN o_sram_wen
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 596.000 101.570 600.000 ;
    END
  END o_sram_wen
  PIN o_wb_dbg_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END o_wb_dbg_ack
  PIN o_wb_dbg_rdt[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 57.840 900.000 58.440 ;
    END
  END o_wb_dbg_rdt[0]
  PIN o_wb_dbg_rdt[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.920 4.000 368.520 ;
    END
  END o_wb_dbg_rdt[10]
  PIN o_wb_dbg_rdt[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.920 4.000 402.520 ;
    END
  END o_wb_dbg_rdt[11]
  PIN o_wb_dbg_rdt[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 0.000 471.870 4.000 ;
    END
  END o_wb_dbg_rdt[12]
  PIN o_wb_dbg_rdt[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 4.000 419.520 ;
    END
  END o_wb_dbg_rdt[13]
  PIN o_wb_dbg_rdt[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 0.000 537.650 4.000 ;
    END
  END o_wb_dbg_rdt[14]
  PIN o_wb_dbg_rdt[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.450 0.000 559.730 4.000 ;
    END
  END o_wb_dbg_rdt[15]
  PIN o_wb_dbg_rdt[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 374.720 900.000 375.320 ;
    END
  END o_wb_dbg_rdt[16]
  PIN o_wb_dbg_rdt[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END o_wb_dbg_rdt[17]
  PIN o_wb_dbg_rdt[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.150 0.000 603.430 4.000 ;
    END
  END o_wb_dbg_rdt[18]
  PIN o_wb_dbg_rdt[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 0.000 647.590 4.000 ;
    END
  END o_wb_dbg_rdt[19]
  PIN o_wb_dbg_rdt[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 91.160 900.000 91.760 ;
    END
  END o_wb_dbg_rdt[1]
  PIN o_wb_dbg_rdt[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 424.360 900.000 424.960 ;
    END
  END o_wb_dbg_rdt[20]
  PIN o_wb_dbg_rdt[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.090 0.000 713.370 4.000 ;
    END
  END o_wb_dbg_rdt[21]
  PIN o_wb_dbg_rdt[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 0.000 757.070 4.000 ;
    END
  END o_wb_dbg_rdt[22]
  PIN o_wb_dbg_rdt[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.280 4.000 539.880 ;
    END
  END o_wb_dbg_rdt[23]
  PIN o_wb_dbg_rdt[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 457.680 900.000 458.280 ;
    END
  END o_wb_dbg_rdt[24]
  PIN o_wb_dbg_rdt[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.280 4.000 556.880 ;
    END
  END o_wb_dbg_rdt[25]
  PIN o_wb_dbg_rdt[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.280 4.000 573.880 ;
    END
  END o_wb_dbg_rdt[26]
  PIN o_wb_dbg_rdt[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 508.000 900.000 508.600 ;
    END
  END o_wb_dbg_rdt[27]
  PIN o_wb_dbg_rdt[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 541.320 900.000 541.920 ;
    END
  END o_wb_dbg_rdt[28]
  PIN o_wb_dbg_rdt[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.150 596.000 856.430 600.000 ;
    END
  END o_wb_dbg_rdt[29]
  PIN o_wb_dbg_rdt[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 596.000 304.890 600.000 ;
    END
  END o_wb_dbg_rdt[2]
  PIN o_wb_dbg_rdt[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 574.640 900.000 575.240 ;
    END
  END o_wb_dbg_rdt[30]
  PIN o_wb_dbg_rdt[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 590.960 900.000 591.560 ;
    END
  END o_wb_dbg_rdt[31]
  PIN o_wb_dbg_rdt[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 174.800 900.000 175.400 ;
    END
  END o_wb_dbg_rdt[3]
  PIN o_wb_dbg_rdt[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END o_wb_dbg_rdt[4]
  PIN o_wb_dbg_rdt[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.870 0.000 296.150 4.000 ;
    END
  END o_wb_dbg_rdt[5]
  PIN o_wb_dbg_rdt[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 596.000 420.810 600.000 ;
    END
  END o_wb_dbg_rdt[6]
  PIN o_wb_dbg_rdt[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 596.000 537.190 600.000 ;
    END
  END o_wb_dbg_rdt[7]
  PIN o_wb_dbg_rdt[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END o_wb_dbg_rdt[8]
  PIN o_wb_dbg_rdt[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END o_wb_dbg_rdt[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 792.340 10.880 793.940 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 638.740 10.880 640.340 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 485.140 10.880 486.740 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.540 10.880 333.140 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 587.520 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 869.140 10.880 870.740 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 715.540 10.880 717.140 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 561.940 10.880 563.540 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 408.340 10.880 409.940 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.740 10.880 256.340 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 587.520 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 795.640 10.880 797.240 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 642.040 10.880 643.640 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 488.440 10.880 490.040 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 334.840 10.880 336.440 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.240 10.880 182.840 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.640 10.880 29.240 587.520 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 872.440 10.880 874.040 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 718.840 10.880 720.440 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 565.240 10.880 566.840 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 411.640 10.880 413.240 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 258.040 10.880 259.640 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.440 10.880 106.040 587.520 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 798.940 10.880 800.540 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 645.340 10.880 646.940 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 491.740 10.880 493.340 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 338.140 10.880 339.740 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.540 10.880 186.140 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.880 32.540 587.520 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 875.740 10.880 877.340 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 722.140 10.880 723.740 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 568.540 10.880 570.140 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 414.940 10.880 416.540 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 261.340 10.880 262.940 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.740 10.880 109.340 587.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 229.225 11.305 885.815 281.775 ;
      LAYER met1 ;
        RECT 5.520 10.640 894.240 587.760 ;
      LAYER met2 ;
        RECT 10.680 595.720 14.070 596.000 ;
        RECT 14.910 595.720 43.050 596.000 ;
        RECT 43.890 595.720 72.030 596.000 ;
        RECT 72.870 595.720 101.010 596.000 ;
        RECT 101.850 595.720 129.990 596.000 ;
        RECT 130.830 595.720 158.970 596.000 ;
        RECT 159.810 595.720 187.950 596.000 ;
        RECT 188.790 595.720 216.930 596.000 ;
        RECT 217.770 595.720 246.370 596.000 ;
        RECT 247.210 595.720 275.350 596.000 ;
        RECT 276.190 595.720 304.330 596.000 ;
        RECT 305.170 595.720 333.310 596.000 ;
        RECT 334.150 595.720 362.290 596.000 ;
        RECT 363.130 595.720 391.270 596.000 ;
        RECT 392.110 595.720 420.250 596.000 ;
        RECT 421.090 595.720 449.230 596.000 ;
        RECT 450.070 595.720 478.670 596.000 ;
        RECT 479.510 595.720 507.650 596.000 ;
        RECT 508.490 595.720 536.630 596.000 ;
        RECT 537.470 595.720 565.610 596.000 ;
        RECT 566.450 595.720 594.590 596.000 ;
        RECT 595.430 595.720 623.570 596.000 ;
        RECT 624.410 595.720 652.550 596.000 ;
        RECT 653.390 595.720 681.530 596.000 ;
        RECT 682.370 595.720 710.970 596.000 ;
        RECT 711.810 595.720 739.950 596.000 ;
        RECT 740.790 595.720 768.930 596.000 ;
        RECT 769.770 595.720 797.910 596.000 ;
        RECT 798.750 595.720 826.890 596.000 ;
        RECT 827.730 595.720 855.870 596.000 ;
        RECT 856.710 595.720 884.850 596.000 ;
        RECT 885.690 595.720 889.020 596.000 ;
        RECT 10.680 4.280 889.020 595.720 ;
        RECT 11.230 4.000 32.010 4.280 ;
        RECT 32.850 4.000 54.090 4.280 ;
        RECT 54.930 4.000 76.170 4.280 ;
        RECT 77.010 4.000 97.790 4.280 ;
        RECT 98.630 4.000 119.870 4.280 ;
        RECT 120.710 4.000 141.950 4.280 ;
        RECT 142.790 4.000 164.030 4.280 ;
        RECT 164.870 4.000 185.650 4.280 ;
        RECT 186.490 4.000 207.730 4.280 ;
        RECT 208.570 4.000 229.810 4.280 ;
        RECT 230.650 4.000 251.890 4.280 ;
        RECT 252.730 4.000 273.510 4.280 ;
        RECT 274.350 4.000 295.590 4.280 ;
        RECT 296.430 4.000 317.670 4.280 ;
        RECT 318.510 4.000 339.290 4.280 ;
        RECT 340.130 4.000 361.370 4.280 ;
        RECT 362.210 4.000 383.450 4.280 ;
        RECT 384.290 4.000 405.530 4.280 ;
        RECT 406.370 4.000 427.150 4.280 ;
        RECT 427.990 4.000 449.230 4.280 ;
        RECT 450.070 4.000 471.310 4.280 ;
        RECT 472.150 4.000 493.390 4.280 ;
        RECT 494.230 4.000 515.010 4.280 ;
        RECT 515.850 4.000 537.090 4.280 ;
        RECT 537.930 4.000 559.170 4.280 ;
        RECT 560.010 4.000 581.250 4.280 ;
        RECT 582.090 4.000 602.870 4.280 ;
        RECT 603.710 4.000 624.950 4.280 ;
        RECT 625.790 4.000 647.030 4.280 ;
        RECT 647.870 4.000 668.650 4.280 ;
        RECT 669.490 4.000 690.730 4.280 ;
        RECT 691.570 4.000 712.810 4.280 ;
        RECT 713.650 4.000 734.890 4.280 ;
        RECT 735.730 4.000 756.510 4.280 ;
        RECT 757.350 4.000 778.590 4.280 ;
        RECT 779.430 4.000 800.670 4.280 ;
        RECT 801.510 4.000 822.750 4.280 ;
        RECT 823.590 4.000 844.370 4.280 ;
        RECT 845.210 4.000 866.450 4.280 ;
        RECT 867.290 4.000 888.530 4.280 ;
      LAYER met3 ;
        RECT 4.000 591.280 895.600 591.425 ;
        RECT 4.400 590.560 895.600 591.280 ;
        RECT 4.400 589.880 896.000 590.560 ;
        RECT 4.000 575.640 896.000 589.880 ;
        RECT 4.000 574.280 895.600 575.640 ;
        RECT 4.400 574.240 895.600 574.280 ;
        RECT 4.400 572.880 896.000 574.240 ;
        RECT 4.000 558.640 896.000 572.880 ;
        RECT 4.000 557.280 895.600 558.640 ;
        RECT 4.400 557.240 895.600 557.280 ;
        RECT 4.400 555.880 896.000 557.240 ;
        RECT 4.000 542.320 896.000 555.880 ;
        RECT 4.000 540.920 895.600 542.320 ;
        RECT 4.000 540.280 896.000 540.920 ;
        RECT 4.400 538.880 896.000 540.280 ;
        RECT 4.000 525.320 896.000 538.880 ;
        RECT 4.000 523.920 895.600 525.320 ;
        RECT 4.000 523.280 896.000 523.920 ;
        RECT 4.400 521.880 896.000 523.280 ;
        RECT 4.000 509.000 896.000 521.880 ;
        RECT 4.000 507.600 895.600 509.000 ;
        RECT 4.000 505.600 896.000 507.600 ;
        RECT 4.400 504.200 896.000 505.600 ;
        RECT 4.000 492.000 896.000 504.200 ;
        RECT 4.000 490.600 895.600 492.000 ;
        RECT 4.000 488.600 896.000 490.600 ;
        RECT 4.400 487.200 896.000 488.600 ;
        RECT 4.000 475.680 896.000 487.200 ;
        RECT 4.000 474.280 895.600 475.680 ;
        RECT 4.000 471.600 896.000 474.280 ;
        RECT 4.400 470.200 896.000 471.600 ;
        RECT 4.000 458.680 896.000 470.200 ;
        RECT 4.000 457.280 895.600 458.680 ;
        RECT 4.000 454.600 896.000 457.280 ;
        RECT 4.400 453.200 896.000 454.600 ;
        RECT 4.000 442.360 896.000 453.200 ;
        RECT 4.000 440.960 895.600 442.360 ;
        RECT 4.000 437.600 896.000 440.960 ;
        RECT 4.400 436.200 896.000 437.600 ;
        RECT 4.000 425.360 896.000 436.200 ;
        RECT 4.000 423.960 895.600 425.360 ;
        RECT 4.000 419.920 896.000 423.960 ;
        RECT 4.400 418.520 896.000 419.920 ;
        RECT 4.000 409.040 896.000 418.520 ;
        RECT 4.000 407.640 895.600 409.040 ;
        RECT 4.000 402.920 896.000 407.640 ;
        RECT 4.400 401.520 896.000 402.920 ;
        RECT 4.000 392.040 896.000 401.520 ;
        RECT 4.000 390.640 895.600 392.040 ;
        RECT 4.000 385.920 896.000 390.640 ;
        RECT 4.400 384.520 896.000 385.920 ;
        RECT 4.000 375.720 896.000 384.520 ;
        RECT 4.000 374.320 895.600 375.720 ;
        RECT 4.000 368.920 896.000 374.320 ;
        RECT 4.400 367.520 896.000 368.920 ;
        RECT 4.000 358.720 896.000 367.520 ;
        RECT 4.000 357.320 895.600 358.720 ;
        RECT 4.000 351.920 896.000 357.320 ;
        RECT 4.400 350.520 896.000 351.920 ;
        RECT 4.000 342.400 896.000 350.520 ;
        RECT 4.000 341.000 895.600 342.400 ;
        RECT 4.000 334.240 896.000 341.000 ;
        RECT 4.400 332.840 896.000 334.240 ;
        RECT 4.000 325.400 896.000 332.840 ;
        RECT 4.000 324.000 895.600 325.400 ;
        RECT 4.000 317.240 896.000 324.000 ;
        RECT 4.400 315.840 896.000 317.240 ;
        RECT 4.000 309.080 896.000 315.840 ;
        RECT 4.000 307.680 895.600 309.080 ;
        RECT 4.000 300.240 896.000 307.680 ;
        RECT 4.400 298.840 896.000 300.240 ;
        RECT 4.000 292.080 896.000 298.840 ;
        RECT 4.000 290.680 895.600 292.080 ;
        RECT 4.000 283.240 896.000 290.680 ;
        RECT 4.400 281.840 896.000 283.240 ;
        RECT 4.000 275.760 896.000 281.840 ;
        RECT 4.000 274.360 895.600 275.760 ;
        RECT 4.000 266.240 896.000 274.360 ;
        RECT 4.400 264.840 896.000 266.240 ;
        RECT 4.000 258.760 896.000 264.840 ;
        RECT 4.000 257.360 895.600 258.760 ;
        RECT 4.000 248.560 896.000 257.360 ;
        RECT 4.400 247.160 896.000 248.560 ;
        RECT 4.000 242.440 896.000 247.160 ;
        RECT 4.000 241.040 895.600 242.440 ;
        RECT 4.000 231.560 896.000 241.040 ;
        RECT 4.400 230.160 896.000 231.560 ;
        RECT 4.000 225.440 896.000 230.160 ;
        RECT 4.000 224.040 895.600 225.440 ;
        RECT 4.000 214.560 896.000 224.040 ;
        RECT 4.400 213.160 896.000 214.560 ;
        RECT 4.000 209.120 896.000 213.160 ;
        RECT 4.000 207.720 895.600 209.120 ;
        RECT 4.000 197.560 896.000 207.720 ;
        RECT 4.400 196.160 896.000 197.560 ;
        RECT 4.000 192.120 896.000 196.160 ;
        RECT 4.000 190.720 895.600 192.120 ;
        RECT 4.000 180.560 896.000 190.720 ;
        RECT 4.400 179.160 896.000 180.560 ;
        RECT 4.000 175.800 896.000 179.160 ;
        RECT 4.000 174.400 895.600 175.800 ;
        RECT 4.000 162.880 896.000 174.400 ;
        RECT 4.400 161.480 896.000 162.880 ;
        RECT 4.000 158.800 896.000 161.480 ;
        RECT 4.000 157.400 895.600 158.800 ;
        RECT 4.000 145.880 896.000 157.400 ;
        RECT 4.400 144.480 896.000 145.880 ;
        RECT 4.000 142.480 896.000 144.480 ;
        RECT 4.000 141.080 895.600 142.480 ;
        RECT 4.000 128.880 896.000 141.080 ;
        RECT 4.400 127.480 896.000 128.880 ;
        RECT 4.000 125.480 896.000 127.480 ;
        RECT 4.000 124.080 895.600 125.480 ;
        RECT 4.000 111.880 896.000 124.080 ;
        RECT 4.400 110.480 896.000 111.880 ;
        RECT 4.000 109.160 896.000 110.480 ;
        RECT 4.000 107.760 895.600 109.160 ;
        RECT 4.000 94.880 896.000 107.760 ;
        RECT 4.400 93.480 896.000 94.880 ;
        RECT 4.000 92.160 896.000 93.480 ;
        RECT 4.000 90.760 895.600 92.160 ;
        RECT 4.000 77.200 896.000 90.760 ;
        RECT 4.400 75.840 896.000 77.200 ;
        RECT 4.400 75.800 895.600 75.840 ;
        RECT 4.000 74.440 895.600 75.800 ;
        RECT 4.000 60.200 896.000 74.440 ;
        RECT 4.400 58.840 896.000 60.200 ;
        RECT 4.400 58.800 895.600 58.840 ;
        RECT 4.000 57.440 895.600 58.800 ;
        RECT 4.000 43.200 896.000 57.440 ;
        RECT 4.400 42.520 896.000 43.200 ;
        RECT 4.400 41.800 895.600 42.520 ;
        RECT 4.000 41.120 895.600 41.800 ;
        RECT 4.000 26.200 896.000 41.120 ;
        RECT 4.400 25.520 896.000 26.200 ;
        RECT 4.400 24.800 895.600 25.520 ;
        RECT 4.000 24.120 895.600 24.800 ;
        RECT 4.000 9.200 896.000 24.120 ;
        RECT 4.400 8.335 895.600 9.200 ;
      LAYER met4 ;
        RECT 46.790 17.175 97.440 579.185 ;
        RECT 99.840 17.175 100.740 579.185 ;
        RECT 103.140 17.175 104.040 579.185 ;
        RECT 106.440 17.175 107.340 579.185 ;
        RECT 109.740 17.175 174.240 579.185 ;
        RECT 176.640 17.175 177.540 579.185 ;
        RECT 179.940 17.175 180.840 579.185 ;
        RECT 183.240 17.175 184.140 579.185 ;
        RECT 186.540 17.175 251.040 579.185 ;
        RECT 253.440 17.175 254.340 579.185 ;
        RECT 256.740 17.175 257.640 579.185 ;
        RECT 260.040 17.175 260.940 579.185 ;
        RECT 263.340 17.175 327.840 579.185 ;
        RECT 330.240 17.175 331.140 579.185 ;
        RECT 333.540 17.175 334.440 579.185 ;
        RECT 336.840 17.175 337.740 579.185 ;
        RECT 340.140 17.175 404.640 579.185 ;
        RECT 407.040 17.175 407.940 579.185 ;
        RECT 410.340 17.175 411.240 579.185 ;
        RECT 413.640 17.175 414.540 579.185 ;
        RECT 416.940 17.175 481.440 579.185 ;
        RECT 483.840 17.175 484.740 579.185 ;
        RECT 487.140 17.175 488.040 579.185 ;
        RECT 490.440 17.175 491.340 579.185 ;
        RECT 493.740 17.175 558.240 579.185 ;
        RECT 560.640 17.175 561.540 579.185 ;
        RECT 563.940 17.175 564.840 579.185 ;
        RECT 567.240 17.175 568.140 579.185 ;
        RECT 570.540 17.175 635.040 579.185 ;
        RECT 637.440 17.175 638.340 579.185 ;
        RECT 640.740 17.175 641.640 579.185 ;
        RECT 644.040 17.175 644.940 579.185 ;
        RECT 647.340 17.175 711.840 579.185 ;
        RECT 714.240 17.175 715.140 579.185 ;
        RECT 717.540 17.175 718.440 579.185 ;
        RECT 720.840 17.175 721.740 579.185 ;
        RECT 724.140 17.175 738.890 579.185 ;
      LAYER met5 ;
        RECT 46.580 235.500 739.100 240.500 ;
  END
END subservient
END LIBRARY

