VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sky130_sram_1kbyte_1rw1r_32x256_8
   CLASS BLOCK ;
   SIZE 462.1 BY 383.22 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  97.92 0.0 98.3 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  104.04 0.0 104.42 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  109.48 0.0 109.86 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  116.28 0.0 116.66 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  121.72 0.0 122.1 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  127.16 0.0 127.54 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  132.6 0.0 132.98 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  139.4 0.0 139.78 0.38 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  144.84 0.0 145.22 0.38 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  150.28 0.0 150.66 0.38 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  156.4 0.0 156.78 0.38 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  161.84 0.0 162.22 0.38 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  168.64 0.0 169.02 0.38 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  174.08 0.0 174.46 0.38 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  179.52 0.0 179.9 0.38 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  185.64 0.0 186.02 0.38 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  192.44 0.0 192.82 0.38 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  197.88 0.0 198.26 0.38 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  203.32 0.0 203.7 0.38 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  208.76 0.0 209.14 0.38 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  215.56 0.0 215.94 0.38 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  221.0 0.0 221.38 0.38 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  226.44 0.0 226.82 0.38 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  232.56 0.0 232.94 0.38 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  238.0 0.0 238.38 0.38 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  244.8 0.0 245.18 0.38 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  250.24 0.0 250.62 0.38 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  255.68 0.0 256.06 0.38 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  261.12 0.0 261.5 0.38 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  267.24 0.0 267.62 0.38 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  274.04 0.0 274.42 0.38 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  279.48 0.0 279.86 0.38 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  68.68 0.0 69.06 0.38 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 121.72 0.38 122.1 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 129.88 0.38 130.26 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 135.32 0.38 135.7 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 143.48 0.38 143.86 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 148.92 0.38 149.3 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 157.76 0.38 158.14 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 163.2 0.38 163.58 ;
      END
   END addr0[7]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  388.28 382.84 388.66 383.22 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  461.72 76.16 462.1 76.54 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  461.72 68.0 462.1 68.38 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  461.72 61.88 462.1 62.26 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  406.64 0.0 407.02 0.38 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  404.6 0.0 404.98 0.38 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  405.28 0.0 405.66 0.38 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  405.96 0.0 406.34 0.38 ;
      END
   END addr1[7]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 21.08 0.38 21.46 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  461.72 375.36 462.1 375.74 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 29.24 0.38 29.62 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  20.4 0.0 20.78 0.38 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  441.32 382.84 441.7 383.22 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  74.8 0.0 75.18 0.38 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  80.24 0.0 80.62 0.38 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  87.04 0.0 87.42 0.38 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  91.8 0.0 92.18 0.38 ;
      END
   END wmask0[3]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  130.56 0.0 130.94 0.38 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  137.36 0.0 137.74 0.38 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  142.8 0.0 143.18 0.38 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  150.96 0.0 151.34 0.38 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  157.08 0.0 157.46 0.38 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  163.2 0.0 163.58 0.38 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  169.32 0.0 169.7 0.38 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  175.44 0.0 175.82 0.38 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  180.2 0.0 180.58 0.38 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  187.68 0.0 188.06 0.38 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  194.48 0.0 194.86 0.38 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  200.6 0.0 200.98 0.38 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  206.72 0.0 207.1 0.38 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  212.84 0.0 213.22 0.38 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  218.96 0.0 219.34 0.38 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  224.4 0.0 224.78 0.38 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  230.52 0.0 230.9 0.38 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  236.64 0.0 237.02 0.38 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  244.12 0.0 244.5 0.38 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  248.2 0.0 248.58 0.38 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  257.04 0.0 257.42 0.38 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  263.16 0.0 263.54 0.38 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  269.28 0.0 269.66 0.38 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  275.4 0.0 275.78 0.38 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  280.16 0.0 280.54 0.38 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  287.64 0.0 288.02 0.38 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  293.76 0.0 294.14 0.38 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  300.56 0.0 300.94 0.38 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  306.68 0.0 307.06 0.38 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  312.8 0.0 313.18 0.38 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  318.92 0.0 319.3 0.38 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  325.04 0.0 325.42 0.38 ;
      END
   END dout0[31]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  131.92 382.84 132.3 383.22 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  138.72 382.84 139.1 383.22 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  144.16 382.84 144.54 383.22 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  150.96 382.84 151.34 383.22 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  157.08 382.84 157.46 383.22 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  163.88 382.84 164.26 383.22 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  170.0 382.84 170.38 383.22 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  175.44 382.84 175.82 383.22 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  182.24 382.84 182.62 383.22 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  187.68 382.84 188.06 383.22 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  194.48 382.84 194.86 383.22 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  200.6 382.84 200.98 383.22 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  207.4 382.84 207.78 383.22 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  212.84 382.84 213.22 383.22 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  218.96 382.84 219.34 383.22 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  225.76 382.84 226.14 383.22 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  231.88 382.84 232.26 383.22 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  238.68 382.84 239.06 383.22 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  244.12 382.84 244.5 383.22 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  250.92 382.84 251.3 383.22 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  256.36 382.84 256.74 383.22 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  262.48 382.84 262.86 383.22 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  269.28 382.84 269.66 383.22 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  275.4 382.84 275.78 383.22 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  282.2 382.84 282.58 383.22 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  287.64 382.84 288.02 383.22 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  294.44 382.84 294.82 383.22 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  300.56 382.84 300.94 383.22 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  307.36 382.84 307.74 383.22 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  312.8 382.84 313.18 383.22 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  318.92 382.84 319.3 383.22 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  325.72 382.84 326.1 383.22 ;
      END
   END dout1[31]
   PIN vcdd1 
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  1.36 0.0 2.42 382.54 ;
      END
   END vcdd1
   PIN vsdd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  0.0 0.0 1.06 382.54 ;
      END
   END vsdd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 461.48 382.6 ;
   LAYER  met2 ;
      RECT  0.62 0.62 461.48 382.6 ;
   LAYER  met3 ;
      RECT  0.68 121.42 461.48 122.4 ;
      RECT  0.62 122.4 0.68 129.58 ;
      RECT  0.62 130.56 0.68 135.02 ;
      RECT  0.62 136.0 0.68 143.18 ;
      RECT  0.62 144.16 0.68 148.62 ;
      RECT  0.62 149.6 0.68 157.46 ;
      RECT  0.62 158.44 0.68 162.9 ;
      RECT  0.62 163.88 0.68 382.6 ;
      RECT  0.68 0.62 461.42 75.86 ;
      RECT  0.68 75.86 461.42 76.84 ;
      RECT  0.68 76.84 461.42 121.42 ;
      RECT  461.42 76.84 461.48 121.42 ;
      RECT  461.42 68.68 461.48 75.86 ;
      RECT  461.42 0.62 461.48 61.58 ;
      RECT  461.42 62.56 461.48 67.7 ;
      RECT  0.62 0.62 0.68 20.78 ;
      RECT  0.68 122.4 461.42 375.06 ;
      RECT  0.68 375.06 461.42 376.04 ;
      RECT  0.68 376.04 461.42 382.6 ;
      RECT  461.42 122.4 461.48 375.06 ;
      RECT  461.42 376.04 461.48 382.6 ;
      RECT  0.62 21.76 0.68 28.94 ;
      RECT  0.62 29.92 0.68 121.42 ;
   LAYER  met4 ;
      RECT  97.62 0.68 98.6 382.6 ;
      RECT  98.6 0.62 103.74 0.68 ;
      RECT  104.72 0.62 109.18 0.68 ;
      RECT  110.16 0.62 115.98 0.68 ;
      RECT  116.96 0.62 121.42 0.68 ;
      RECT  122.4 0.62 126.86 0.68 ;
      RECT  145.52 0.62 149.98 0.68 ;
      RECT  250.92 0.62 255.38 0.68 ;
      RECT  98.6 0.68 387.98 382.54 ;
      RECT  387.98 0.68 388.96 382.54 ;
      RECT  388.96 0.68 461.48 382.54 ;
      RECT  407.32 0.62 461.48 0.68 ;
      RECT  21.08 0.62 68.38 0.68 ;
      RECT  388.96 382.54 441.02 382.6 ;
      RECT  442.0 382.54 461.48 382.6 ;
      RECT  69.36 0.62 74.5 0.68 ;
      RECT  75.48 0.62 79.94 0.68 ;
      RECT  80.92 0.62 86.74 0.68 ;
      RECT  87.72 0.62 91.5 0.68 ;
      RECT  92.48 0.62 97.62 0.68 ;
      RECT  127.84 0.62 130.26 0.68 ;
      RECT  131.24 0.62 132.3 0.68 ;
      RECT  133.28 0.62 137.06 0.68 ;
      RECT  138.04 0.62 139.1 0.68 ;
      RECT  140.08 0.62 142.5 0.68 ;
      RECT  143.48 0.62 144.54 0.68 ;
      RECT  151.64 0.62 156.1 0.68 ;
      RECT  157.76 0.62 161.54 0.68 ;
      RECT  162.52 0.62 162.9 0.68 ;
      RECT  163.88 0.62 168.34 0.68 ;
      RECT  170.0 0.62 173.78 0.68 ;
      RECT  174.76 0.62 175.14 0.68 ;
      RECT  176.12 0.62 179.22 0.68 ;
      RECT  180.88 0.62 185.34 0.68 ;
      RECT  186.32 0.62 187.38 0.68 ;
      RECT  188.36 0.62 192.14 0.68 ;
      RECT  193.12 0.62 194.18 0.68 ;
      RECT  195.16 0.62 197.58 0.68 ;
      RECT  198.56 0.62 200.3 0.68 ;
      RECT  201.28 0.62 203.02 0.68 ;
      RECT  204.0 0.62 206.42 0.68 ;
      RECT  207.4 0.62 208.46 0.68 ;
      RECT  209.44 0.62 212.54 0.68 ;
      RECT  213.52 0.62 215.26 0.68 ;
      RECT  216.24 0.62 218.66 0.68 ;
      RECT  219.64 0.62 220.7 0.68 ;
      RECT  221.68 0.62 224.1 0.68 ;
      RECT  225.08 0.62 226.14 0.68 ;
      RECT  227.12 0.62 230.22 0.68 ;
      RECT  231.2 0.62 232.26 0.68 ;
      RECT  233.24 0.62 236.34 0.68 ;
      RECT  237.32 0.62 237.7 0.68 ;
      RECT  238.68 0.62 243.82 0.68 ;
      RECT  245.48 0.62 247.9 0.68 ;
      RECT  248.88 0.62 249.94 0.68 ;
      RECT  256.36 0.62 256.74 0.68 ;
      RECT  257.72 0.62 260.82 0.68 ;
      RECT  261.8 0.62 262.86 0.68 ;
      RECT  263.84 0.62 266.94 0.68 ;
      RECT  267.92 0.62 268.98 0.68 ;
      RECT  269.96 0.62 273.74 0.68 ;
      RECT  274.72 0.62 275.1 0.68 ;
      RECT  276.08 0.62 279.18 0.68 ;
      RECT  280.84 0.62 287.34 0.68 ;
      RECT  288.32 0.62 293.46 0.68 ;
      RECT  294.44 0.62 300.26 0.68 ;
      RECT  301.24 0.62 306.38 0.68 ;
      RECT  307.36 0.62 312.5 0.68 ;
      RECT  313.48 0.62 318.62 0.68 ;
      RECT  319.6 0.62 324.74 0.68 ;
      RECT  325.72 0.62 404.3 0.68 ;
      RECT  98.6 382.54 131.62 382.6 ;
      RECT  132.6 382.54 138.42 382.6 ;
      RECT  139.4 382.54 143.86 382.6 ;
      RECT  144.84 382.54 150.66 382.6 ;
      RECT  151.64 382.54 156.78 382.6 ;
      RECT  157.76 382.54 163.58 382.6 ;
      RECT  164.56 382.54 169.7 382.6 ;
      RECT  170.68 382.54 175.14 382.6 ;
      RECT  176.12 382.54 181.94 382.6 ;
      RECT  182.92 382.54 187.38 382.6 ;
      RECT  188.36 382.54 194.18 382.6 ;
      RECT  195.16 382.54 200.3 382.6 ;
      RECT  201.28 382.54 207.1 382.6 ;
      RECT  208.08 382.54 212.54 382.6 ;
      RECT  213.52 382.54 218.66 382.6 ;
      RECT  219.64 382.54 225.46 382.6 ;
      RECT  226.44 382.54 231.58 382.6 ;
      RECT  232.56 382.54 238.38 382.6 ;
      RECT  239.36 382.54 243.82 382.6 ;
      RECT  244.8 382.54 250.62 382.6 ;
      RECT  251.6 382.54 256.06 382.6 ;
      RECT  257.04 382.54 262.18 382.6 ;
      RECT  263.16 382.54 268.98 382.6 ;
      RECT  269.96 382.54 275.1 382.6 ;
      RECT  276.08 382.54 281.9 382.6 ;
      RECT  282.88 382.54 287.34 382.6 ;
      RECT  288.32 382.54 294.14 382.6 ;
      RECT  295.12 382.54 300.26 382.6 ;
      RECT  301.24 382.54 307.06 382.6 ;
      RECT  308.04 382.54 312.5 382.6 ;
      RECT  313.48 382.54 318.62 382.6 ;
      RECT  319.6 382.54 325.42 382.6 ;
      RECT  326.4 382.54 387.98 382.6 ;
      RECT  2.72 0.68 97.62 382.6 ;
      RECT  2.72 0.62 20.1 0.68 ;
   END
END    sky130_sram_1kbyte_1rw1r_32x256_8
END    LIBRARY
