VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO subservient
  CLASS BLOCK ;
  FOREIGN subservient ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN i_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 596.000 10.490 600.000 ;
    END
  END i_clk
  PIN i_debug_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 4.000 ;
    END
  END i_debug_mode
  PIN i_dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 6.840 900.000 7.440 ;
    END
  END i_dout1[0]
  PIN i_dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 306.720 900.000 307.320 ;
    END
  END i_dout1[10]
  PIN i_dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 321.000 900.000 321.600 ;
    END
  END i_dout1[11]
  PIN i_dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 0.000 465.890 4.000 ;
    END
  END i_dout1[12]
  PIN i_dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END i_dout1[13]
  PIN i_dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 596.000 419.430 600.000 ;
    END
  END i_dout1[14]
  PIN i_dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 305.360 4.000 305.960 ;
    END
  END i_dout1[15]
  PIN i_dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.330 596.000 480.610 600.000 ;
    END
  END i_dout1[16]
  PIN i_dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.970 596.000 542.250 600.000 ;
    END
  END i_dout1[17]
  PIN i_dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 0.000 592.390 4.000 ;
    END
  END i_dout1[18]
  PIN i_dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 392.400 900.000 393.000 ;
    END
  END i_dout1[19]
  PIN i_dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 21.120 900.000 21.720 ;
    END
  END i_dout1[1]
  PIN i_dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END i_dout1[20]
  PIN i_dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.800 4.000 413.400 ;
    END
  END i_dout1[21]
  PIN i_dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.280 4.000 437.880 ;
    END
  END i_dout1[22]
  PIN i_dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.970 596.000 726.250 600.000 ;
    END
  END i_dout1[23]
  PIN i_dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 449.520 900.000 450.120 ;
    END
  END i_dout1[24]
  PIN i_dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.080 4.000 461.680 ;
    END
  END i_dout1[25]
  PIN i_dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.880 4.000 485.480 ;
    END
  END i_dout1[26]
  PIN i_dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.160 4.000 533.760 ;
    END
  END i_dout1[27]
  PIN i_dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.720 4.000 545.320 ;
    END
  END i_dout1[28]
  PIN i_dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.390 0.000 876.670 4.000 ;
    END
  END i_dout1[29]
  PIN i_dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 35.400 900.000 36.000 ;
    END
  END i_dout1[2]
  PIN i_dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.790 596.000 849.070 600.000 ;
    END
  END i_dout1[30]
  PIN i_dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 578.040 900.000 578.640 ;
    END
  END i_dout1[31]
  PIN i_dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 49.680 900.000 50.280 ;
    END
  END i_dout1[3]
  PIN i_dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END i_dout1[4]
  PIN i_dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END i_dout1[5]
  PIN i_dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END i_dout1[6]
  PIN i_dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END i_dout1[7]
  PIN i_dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 596.000 337.550 600.000 ;
    END
  END i_dout1[8]
  PIN i_dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END i_dout1[9]
  PIN i_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 4.000 ;
    END
  END i_rst
  PIN i_wb_dbg_adr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END i_wb_dbg_adr[0]
  PIN i_wb_dbg_adr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END i_wb_dbg_adr[10]
  PIN i_wb_dbg_adr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 0.000 434.610 4.000 ;
    END
  END i_wb_dbg_adr[11]
  PIN i_wb_dbg_adr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 0.000 481.990 4.000 ;
    END
  END i_wb_dbg_adr[12]
  PIN i_wb_dbg_adr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 349.560 900.000 350.160 ;
    END
  END i_wb_dbg_adr[13]
  PIN i_wb_dbg_adr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 363.840 900.000 364.440 ;
    END
  END i_wb_dbg_adr[14]
  PIN i_wb_dbg_adr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 596.000 460.370 600.000 ;
    END
  END i_wb_dbg_adr[15]
  PIN i_wb_dbg_adr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.030 596.000 501.310 600.000 ;
    END
  END i_wb_dbg_adr[16]
  PIN i_wb_dbg_adr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.960 4.000 353.560 ;
    END
  END i_wb_dbg_adr[17]
  PIN i_wb_dbg_adr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.750 0.000 608.030 4.000 ;
    END
  END i_wb_dbg_adr[18]
  PIN i_wb_dbg_adr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.490 0.000 639.770 4.000 ;
    END
  END i_wb_dbg_adr[19]
  PIN i_wb_dbg_adr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 78.240 900.000 78.840 ;
    END
  END i_wb_dbg_adr[1]
  PIN i_wb_dbg_adr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 406.680 900.000 407.280 ;
    END
  END i_wb_dbg_adr[20]
  PIN i_wb_dbg_adr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 420.960 900.000 421.560 ;
    END
  END i_wb_dbg_adr[21]
  PIN i_wb_dbg_adr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.790 596.000 665.070 600.000 ;
    END
  END i_wb_dbg_adr[22]
  PIN i_wb_dbg_adr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.670 596.000 746.950 600.000 ;
    END
  END i_wb_dbg_adr[23]
  PIN i_wb_dbg_adr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.910 596.000 767.190 600.000 ;
    END
  END i_wb_dbg_adr[24]
  PIN i_wb_dbg_adr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 478.080 900.000 478.680 ;
    END
  END i_wb_dbg_adr[25]
  PIN i_wb_dbg_adr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.850 596.000 808.130 600.000 ;
    END
  END i_wb_dbg_adr[26]
  PIN i_wb_dbg_adr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.270 0.000 797.550 4.000 ;
    END
  END i_wb_dbg_adr[27]
  PIN i_wb_dbg_adr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.960 4.000 557.560 ;
    END
  END i_wb_dbg_adr[28]
  PIN i_wb_dbg_adr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 0.000 892.310 4.000 ;
    END
  END i_wb_dbg_adr[29]
  PIN i_wb_dbg_adr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 106.800 900.000 107.400 ;
    END
  END i_wb_dbg_adr[2]
  PIN i_wb_dbg_adr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 596.000 869.770 600.000 ;
    END
  END i_wb_dbg_adr[30]
  PIN i_wb_dbg_adr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 592.320 900.000 592.920 ;
    END
  END i_wb_dbg_adr[31]
  PIN i_wb_dbg_adr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 596.000 173.790 600.000 ;
    END
  END i_wb_dbg_adr[3]
  PIN i_wb_dbg_adr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END i_wb_dbg_adr[4]
  PIN i_wb_dbg_adr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.200 4.000 161.800 ;
    END
  END i_wb_dbg_adr[5]
  PIN i_wb_dbg_adr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END i_wb_dbg_adr[6]
  PIN i_wb_dbg_adr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 596.000 255.670 600.000 ;
    END
  END i_wb_dbg_adr[7]
  PIN i_wb_dbg_adr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 4.000 ;
    END
  END i_wb_dbg_adr[8]
  PIN i_wb_dbg_adr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 292.440 900.000 293.040 ;
    END
  END i_wb_dbg_adr[9]
  PIN i_wb_dbg_dat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 63.960 900.000 64.560 ;
    END
  END i_wb_dbg_dat[0]
  PIN i_wb_dbg_dat[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 0.000 418.510 4.000 ;
    END
  END i_wb_dbg_dat[10]
  PIN i_wb_dbg_dat[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END i_wb_dbg_dat[11]
  PIN i_wb_dbg_dat[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 0.000 497.630 4.000 ;
    END
  END i_wb_dbg_dat[12]
  PIN i_wb_dbg_dat[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 0.000 513.270 4.000 ;
    END
  END i_wb_dbg_dat[13]
  PIN i_wb_dbg_dat[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.090 0.000 529.370 4.000 ;
    END
  END i_wb_dbg_dat[14]
  PIN i_wb_dbg_dat[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END i_wb_dbg_dat[15]
  PIN i_wb_dbg_dat[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 596.000 521.550 600.000 ;
    END
  END i_wb_dbg_dat[16]
  PIN i_wb_dbg_dat[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 0.000 576.750 4.000 ;
    END
  END i_wb_dbg_dat[17]
  PIN i_wb_dbg_dat[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 596.000 583.190 600.000 ;
    END
  END i_wb_dbg_dat[18]
  PIN i_wb_dbg_dat[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.130 0.000 655.410 4.000 ;
    END
  END i_wb_dbg_dat[19]
  PIN i_wb_dbg_dat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 4.000 ;
    END
  END i_wb_dbg_dat[1]
  PIN i_wb_dbg_dat[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END i_wb_dbg_dat[20]
  PIN i_wb_dbg_dat[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 435.240 900.000 435.840 ;
    END
  END i_wb_dbg_dat[21]
  PIN i_wb_dbg_dat[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 596.000 685.310 600.000 ;
    END
  END i_wb_dbg_dat[22]
  PIN i_wb_dbg_dat[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.610 0.000 718.890 4.000 ;
    END
  END i_wb_dbg_dat[23]
  PIN i_wb_dbg_dat[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 463.800 900.000 464.400 ;
    END
  END i_wb_dbg_dat[24]
  PIN i_wb_dbg_dat[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 0.000 766.270 4.000 ;
    END
  END i_wb_dbg_dat[25]
  PIN i_wb_dbg_dat[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.120 4.000 497.720 ;
    END
  END i_wb_dbg_dat[26]
  PIN i_wb_dbg_dat[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 492.360 900.000 492.960 ;
    END
  END i_wb_dbg_dat[27]
  PIN i_wb_dbg_dat[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.200 4.000 569.800 ;
    END
  END i_wb_dbg_dat[28]
  PIN i_wb_dbg_dat[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 506.640 900.000 507.240 ;
    END
  END i_wb_dbg_dat[29]
  PIN i_wb_dbg_dat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END i_wb_dbg_dat[2]
  PIN i_wb_dbg_dat[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 535.200 900.000 535.800 ;
    END
  END i_wb_dbg_dat[30]
  PIN i_wb_dbg_dat[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 580.760 4.000 581.360 ;
    END
  END i_wb_dbg_dat[31]
  PIN i_wb_dbg_dat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END i_wb_dbg_dat[3]
  PIN i_wb_dbg_dat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END i_wb_dbg_dat[4]
  PIN i_wb_dbg_dat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 192.480 900.000 193.080 ;
    END
  END i_wb_dbg_dat[5]
  PIN i_wb_dbg_dat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 221.040 900.000 221.640 ;
    END
  END i_wb_dbg_dat[6]
  PIN i_wb_dbg_dat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END i_wb_dbg_dat[7]
  PIN i_wb_dbg_dat[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 0.000 355.490 4.000 ;
    END
  END i_wb_dbg_dat[8]
  PIN i_wb_dbg_dat[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 0.000 371.130 4.000 ;
    END
  END i_wb_dbg_dat[9]
  PIN i_wb_dbg_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 596.000 50.970 600.000 ;
    END
  END i_wb_dbg_sel[0]
  PIN i_wb_dbg_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 596.000 91.910 600.000 ;
    END
  END i_wb_dbg_sel[1]
  PIN i_wb_dbg_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 596.000 112.610 600.000 ;
    END
  END i_wb_dbg_sel[2]
  PIN i_wb_dbg_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 149.640 900.000 150.240 ;
    END
  END i_wb_dbg_sel[3]
  PIN i_wb_dbg_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END i_wb_dbg_stb
  PIN i_wb_dbg_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END i_wb_dbg_we
  PIN o_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END o_addr1[0]
  PIN o_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 4.000 ;
    END
  END o_addr1[1]
  PIN o_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 121.080 900.000 121.680 ;
    END
  END o_addr1[2]
  PIN o_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 596.000 194.490 600.000 ;
    END
  END o_addr1[3]
  PIN o_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 178.200 900.000 178.800 ;
    END
  END o_addr1[4]
  PIN o_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 206.760 900.000 207.360 ;
    END
  END o_addr1[5]
  PIN o_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 235.320 900.000 235.920 ;
    END
  END o_addr1[6]
  PIN o_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 596.000 276.370 600.000 ;
    END
  END o_addr1[7]
  PIN o_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END o_csb0
  PIN o_csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END o_csb1
  PIN o_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END o_din0[0]
  PIN o_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.280 4.000 233.880 ;
    END
  END o_din0[10]
  PIN o_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 0.000 450.250 4.000 ;
    END
  END o_din0[11]
  PIN o_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.880 4.000 281.480 ;
    END
  END o_din0[12]
  PIN o_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 596.000 378.490 600.000 ;
    END
  END o_din0[13]
  PIN o_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 596.000 440.130 600.000 ;
    END
  END o_din0[14]
  PIN o_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END o_din0[15]
  PIN o_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.720 4.000 341.320 ;
    END
  END o_din0[16]
  PIN o_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.200 4.000 365.800 ;
    END
  END o_din0[17]
  PIN o_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END o_din0[18]
  PIN o_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.150 596.000 603.430 600.000 ;
    END
  END o_din0[19]
  PIN o_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END o_din0[1]
  PIN o_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 596.000 624.130 600.000 ;
    END
  END o_din0[20]
  PIN o_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 596.000 644.370 600.000 ;
    END
  END o_din0[21]
  PIN o_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 0.000 702.790 4.000 ;
    END
  END o_din0[22]
  PIN o_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 4.000 ;
    END
  END o_din0[23]
  PIN o_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.610 596.000 787.890 600.000 ;
    END
  END o_din0[24]
  PIN o_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END o_din0[25]
  PIN o_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.680 4.000 509.280 ;
    END
  END o_din0[26]
  PIN o_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.370 0.000 813.650 4.000 ;
    END
  END o_din0[27]
  PIN o_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.650 0.000 844.930 4.000 ;
    END
  END o_din0[28]
  PIN o_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.550 596.000 828.830 600.000 ;
    END
  END o_din0[29]
  PIN o_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 596.000 132.850 600.000 ;
    END
  END o_din0[2]
  PIN o_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 549.480 900.000 550.080 ;
    END
  END o_din0[30]
  PIN o_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 593.000 4.000 593.600 ;
    END
  END o_din0[31]
  PIN o_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 4.000 ;
    END
  END o_din0[3]
  PIN o_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END o_din0[4]
  PIN o_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END o_din0[5]
  PIN o_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 0.000 308.110 4.000 ;
    END
  END o_din0[6]
  PIN o_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 596.000 296.610 600.000 ;
    END
  END o_din0[7]
  PIN o_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 278.160 900.000 278.760 ;
    END
  END o_din0[8]
  PIN o_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 596.000 358.250 600.000 ;
    END
  END o_din0[9]
  PIN o_gpio
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 596.000 30.730 600.000 ;
    END
  END o_gpio
  PIN o_waddr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 596.000 71.670 600.000 ;
    END
  END o_waddr0[0]
  PIN o_waddr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END o_waddr0[1]
  PIN o_waddr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 135.360 900.000 135.960 ;
    END
  END o_waddr0[2]
  PIN o_waddr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 4.000 ;
    END
  END o_waddr0[3]
  PIN o_waddr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 596.000 214.730 600.000 ;
    END
  END o_waddr0[4]
  PIN o_waddr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 4.000 ;
    END
  END o_waddr0[5]
  PIN o_waddr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 249.600 900.000 250.200 ;
    END
  END o_waddr0[6]
  PIN o_waddr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 596.000 317.310 600.000 ;
    END
  END o_waddr0[7]
  PIN o_wb_dbg_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END o_wb_dbg_ack
  PIN o_wb_dbg_rdt[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END o_wb_dbg_rdt[0]
  PIN o_wb_dbg_rdt[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END o_wb_dbg_rdt[10]
  PIN o_wb_dbg_rdt[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END o_wb_dbg_rdt[11]
  PIN o_wb_dbg_rdt[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 335.280 900.000 335.880 ;
    END
  END o_wb_dbg_rdt[12]
  PIN o_wb_dbg_rdt[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 596.000 399.190 600.000 ;
    END
  END o_wb_dbg_rdt[13]
  PIN o_wb_dbg_rdt[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.730 0.000 545.010 4.000 ;
    END
  END o_wb_dbg_rdt[14]
  PIN o_wb_dbg_rdt[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END o_wb_dbg_rdt[15]
  PIN o_wb_dbg_rdt[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 378.120 900.000 378.720 ;
    END
  END o_wb_dbg_rdt[16]
  PIN o_wb_dbg_rdt[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.210 596.000 562.490 600.000 ;
    END
  END o_wb_dbg_rdt[17]
  PIN o_wb_dbg_rdt[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 0.000 624.130 4.000 ;
    END
  END o_wb_dbg_rdt[18]
  PIN o_wb_dbg_rdt[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.230 0.000 671.510 4.000 ;
    END
  END o_wb_dbg_rdt[19]
  PIN o_wb_dbg_rdt[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END o_wb_dbg_rdt[1]
  PIN o_wb_dbg_rdt[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.870 0.000 687.150 4.000 ;
    END
  END o_wb_dbg_rdt[20]
  PIN o_wb_dbg_rdt[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END o_wb_dbg_rdt[21]
  PIN o_wb_dbg_rdt[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.730 596.000 706.010 600.000 ;
    END
  END o_wb_dbg_rdt[22]
  PIN o_wb_dbg_rdt[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END o_wb_dbg_rdt[23]
  PIN o_wb_dbg_rdt[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 0.000 750.170 4.000 ;
    END
  END o_wb_dbg_rdt[24]
  PIN o_wb_dbg_rdt[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.630 0.000 781.910 4.000 ;
    END
  END o_wb_dbg_rdt[25]
  PIN o_wb_dbg_rdt[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.920 4.000 521.520 ;
    END
  END o_wb_dbg_rdt[26]
  PIN o_wb_dbg_rdt[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.010 0.000 829.290 4.000 ;
    END
  END o_wb_dbg_rdt[27]
  PIN o_wb_dbg_rdt[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.750 0.000 861.030 4.000 ;
    END
  END o_wb_dbg_rdt[28]
  PIN o_wb_dbg_rdt[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 520.920 900.000 521.520 ;
    END
  END o_wb_dbg_rdt[29]
  PIN o_wb_dbg_rdt[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END o_wb_dbg_rdt[2]
  PIN o_wb_dbg_rdt[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 563.760 900.000 564.360 ;
    END
  END o_wb_dbg_rdt[30]
  PIN o_wb_dbg_rdt[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.730 596.000 890.010 600.000 ;
    END
  END o_wb_dbg_rdt[31]
  PIN o_wb_dbg_rdt[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 163.920 900.000 164.520 ;
    END
  END o_wb_dbg_rdt[3]
  PIN o_wb_dbg_rdt[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 596.000 235.430 600.000 ;
    END
  END o_wb_dbg_rdt[4]
  PIN o_wb_dbg_rdt[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END o_wb_dbg_rdt[5]
  PIN o_wb_dbg_rdt[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 0.000 323.750 4.000 ;
    END
  END o_wb_dbg_rdt[6]
  PIN o_wb_dbg_rdt[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 263.880 900.000 264.480 ;
    END
  END o_wb_dbg_rdt[7]
  PIN o_wb_dbg_rdt[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.800 4.000 209.400 ;
    END
  END o_wb_dbg_rdt[8]
  PIN o_wb_dbg_rdt[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 0.000 387.230 4.000 ;
    END
  END o_wb_dbg_rdt[9]
  PIN o_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END o_wmask0[0]
  PIN o_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 92.520 900.000 93.120 ;
    END
  END o_wmask0[1]
  PIN o_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 596.000 153.550 600.000 ;
    END
  END o_wmask0[2]
  PIN o_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END o_wmask0[3]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 792.340 10.880 793.940 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 638.740 10.880 640.340 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 485.140 10.880 486.740 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.540 10.880 333.140 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 587.520 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 869.140 10.880 870.740 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 715.540 10.880 717.140 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 561.940 10.880 563.540 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 408.340 10.880 409.940 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.740 10.880 256.340 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 587.520 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 795.640 10.880 797.240 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 642.040 10.880 643.640 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 488.440 10.880 490.040 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 334.840 10.880 336.440 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.240 10.880 182.840 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.640 10.880 29.240 587.520 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 872.440 10.880 874.040 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 718.840 10.880 720.440 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 565.240 10.880 566.840 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 411.640 10.880 413.240 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 258.040 10.880 259.640 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.440 10.880 106.040 587.520 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 798.940 10.880 800.540 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 645.340 10.880 646.940 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 491.740 10.880 493.340 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 338.140 10.880 339.740 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.540 10.880 186.140 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.880 32.540 587.520 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 875.740 10.880 877.340 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 722.140 10.880 723.740 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 568.540 10.880 570.140 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 414.940 10.880 416.540 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 261.340 10.880 262.940 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.740 10.880 109.340 587.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 894.240 587.605 ;
      LAYER met1 ;
        RECT 5.520 10.640 894.240 587.760 ;
      LAYER met2 ;
        RECT 7.920 595.720 9.930 596.000 ;
        RECT 10.770 595.720 30.170 596.000 ;
        RECT 31.010 595.720 50.410 596.000 ;
        RECT 51.250 595.720 71.110 596.000 ;
        RECT 71.950 595.720 91.350 596.000 ;
        RECT 92.190 595.720 112.050 596.000 ;
        RECT 112.890 595.720 132.290 596.000 ;
        RECT 133.130 595.720 152.990 596.000 ;
        RECT 153.830 595.720 173.230 596.000 ;
        RECT 174.070 595.720 193.930 596.000 ;
        RECT 194.770 595.720 214.170 596.000 ;
        RECT 215.010 595.720 234.870 596.000 ;
        RECT 235.710 595.720 255.110 596.000 ;
        RECT 255.950 595.720 275.810 596.000 ;
        RECT 276.650 595.720 296.050 596.000 ;
        RECT 296.890 595.720 316.750 596.000 ;
        RECT 317.590 595.720 336.990 596.000 ;
        RECT 337.830 595.720 357.690 596.000 ;
        RECT 358.530 595.720 377.930 596.000 ;
        RECT 378.770 595.720 398.630 596.000 ;
        RECT 399.470 595.720 418.870 596.000 ;
        RECT 419.710 595.720 439.570 596.000 ;
        RECT 440.410 595.720 459.810 596.000 ;
        RECT 460.650 595.720 480.050 596.000 ;
        RECT 480.890 595.720 500.750 596.000 ;
        RECT 501.590 595.720 520.990 596.000 ;
        RECT 521.830 595.720 541.690 596.000 ;
        RECT 542.530 595.720 561.930 596.000 ;
        RECT 562.770 595.720 582.630 596.000 ;
        RECT 583.470 595.720 602.870 596.000 ;
        RECT 603.710 595.720 623.570 596.000 ;
        RECT 624.410 595.720 643.810 596.000 ;
        RECT 644.650 595.720 664.510 596.000 ;
        RECT 665.350 595.720 684.750 596.000 ;
        RECT 685.590 595.720 705.450 596.000 ;
        RECT 706.290 595.720 725.690 596.000 ;
        RECT 726.530 595.720 746.390 596.000 ;
        RECT 747.230 595.720 766.630 596.000 ;
        RECT 767.470 595.720 787.330 596.000 ;
        RECT 788.170 595.720 807.570 596.000 ;
        RECT 808.410 595.720 828.270 596.000 ;
        RECT 829.110 595.720 848.510 596.000 ;
        RECT 849.350 595.720 869.210 596.000 ;
        RECT 870.050 595.720 889.450 596.000 ;
        RECT 7.920 4.280 890.000 595.720 ;
        RECT 8.470 4.000 23.270 4.280 ;
        RECT 24.110 4.000 38.910 4.280 ;
        RECT 39.750 4.000 55.010 4.280 ;
        RECT 55.850 4.000 70.650 4.280 ;
        RECT 71.490 4.000 86.290 4.280 ;
        RECT 87.130 4.000 102.390 4.280 ;
        RECT 103.230 4.000 118.030 4.280 ;
        RECT 118.870 4.000 133.670 4.280 ;
        RECT 134.510 4.000 149.770 4.280 ;
        RECT 150.610 4.000 165.410 4.280 ;
        RECT 166.250 4.000 181.050 4.280 ;
        RECT 181.890 4.000 197.150 4.280 ;
        RECT 197.990 4.000 212.790 4.280 ;
        RECT 213.630 4.000 228.430 4.280 ;
        RECT 229.270 4.000 244.530 4.280 ;
        RECT 245.370 4.000 260.170 4.280 ;
        RECT 261.010 4.000 275.810 4.280 ;
        RECT 276.650 4.000 291.910 4.280 ;
        RECT 292.750 4.000 307.550 4.280 ;
        RECT 308.390 4.000 323.190 4.280 ;
        RECT 324.030 4.000 339.290 4.280 ;
        RECT 340.130 4.000 354.930 4.280 ;
        RECT 355.770 4.000 370.570 4.280 ;
        RECT 371.410 4.000 386.670 4.280 ;
        RECT 387.510 4.000 402.310 4.280 ;
        RECT 403.150 4.000 417.950 4.280 ;
        RECT 418.790 4.000 434.050 4.280 ;
        RECT 434.890 4.000 449.690 4.280 ;
        RECT 450.530 4.000 465.330 4.280 ;
        RECT 466.170 4.000 481.430 4.280 ;
        RECT 482.270 4.000 497.070 4.280 ;
        RECT 497.910 4.000 512.710 4.280 ;
        RECT 513.550 4.000 528.810 4.280 ;
        RECT 529.650 4.000 544.450 4.280 ;
        RECT 545.290 4.000 560.090 4.280 ;
        RECT 560.930 4.000 576.190 4.280 ;
        RECT 577.030 4.000 591.830 4.280 ;
        RECT 592.670 4.000 607.470 4.280 ;
        RECT 608.310 4.000 623.570 4.280 ;
        RECT 624.410 4.000 639.210 4.280 ;
        RECT 640.050 4.000 654.850 4.280 ;
        RECT 655.690 4.000 670.950 4.280 ;
        RECT 671.790 4.000 686.590 4.280 ;
        RECT 687.430 4.000 702.230 4.280 ;
        RECT 703.070 4.000 718.330 4.280 ;
        RECT 719.170 4.000 733.970 4.280 ;
        RECT 734.810 4.000 749.610 4.280 ;
        RECT 750.450 4.000 765.710 4.280 ;
        RECT 766.550 4.000 781.350 4.280 ;
        RECT 782.190 4.000 796.990 4.280 ;
        RECT 797.830 4.000 813.090 4.280 ;
        RECT 813.930 4.000 828.730 4.280 ;
        RECT 829.570 4.000 844.370 4.280 ;
        RECT 845.210 4.000 860.470 4.280 ;
        RECT 861.310 4.000 876.110 4.280 ;
        RECT 876.950 4.000 890.000 4.280 ;
      LAYER met3 ;
        RECT 4.400 593.320 896.000 593.465 ;
        RECT 4.400 592.600 895.600 593.320 ;
        RECT 4.000 591.920 895.600 592.600 ;
        RECT 4.000 581.760 896.000 591.920 ;
        RECT 4.400 580.360 896.000 581.760 ;
        RECT 4.000 579.040 896.000 580.360 ;
        RECT 4.000 577.640 895.600 579.040 ;
        RECT 4.000 570.200 896.000 577.640 ;
        RECT 4.400 568.800 896.000 570.200 ;
        RECT 4.000 564.760 896.000 568.800 ;
        RECT 4.000 563.360 895.600 564.760 ;
        RECT 4.000 557.960 896.000 563.360 ;
        RECT 4.400 556.560 896.000 557.960 ;
        RECT 4.000 550.480 896.000 556.560 ;
        RECT 4.000 549.080 895.600 550.480 ;
        RECT 4.000 545.720 896.000 549.080 ;
        RECT 4.400 544.320 896.000 545.720 ;
        RECT 4.000 536.200 896.000 544.320 ;
        RECT 4.000 534.800 895.600 536.200 ;
        RECT 4.000 534.160 896.000 534.800 ;
        RECT 4.400 532.760 896.000 534.160 ;
        RECT 4.000 521.920 896.000 532.760 ;
        RECT 4.400 520.520 895.600 521.920 ;
        RECT 4.000 509.680 896.000 520.520 ;
        RECT 4.400 508.280 896.000 509.680 ;
        RECT 4.000 507.640 896.000 508.280 ;
        RECT 4.000 506.240 895.600 507.640 ;
        RECT 4.000 498.120 896.000 506.240 ;
        RECT 4.400 496.720 896.000 498.120 ;
        RECT 4.000 493.360 896.000 496.720 ;
        RECT 4.000 491.960 895.600 493.360 ;
        RECT 4.000 485.880 896.000 491.960 ;
        RECT 4.400 484.480 896.000 485.880 ;
        RECT 4.000 479.080 896.000 484.480 ;
        RECT 4.000 477.680 895.600 479.080 ;
        RECT 4.000 473.640 896.000 477.680 ;
        RECT 4.400 472.240 896.000 473.640 ;
        RECT 4.000 464.800 896.000 472.240 ;
        RECT 4.000 463.400 895.600 464.800 ;
        RECT 4.000 462.080 896.000 463.400 ;
        RECT 4.400 460.680 896.000 462.080 ;
        RECT 4.000 450.520 896.000 460.680 ;
        RECT 4.000 449.840 895.600 450.520 ;
        RECT 4.400 449.120 895.600 449.840 ;
        RECT 4.400 448.440 896.000 449.120 ;
        RECT 4.000 438.280 896.000 448.440 ;
        RECT 4.400 436.880 896.000 438.280 ;
        RECT 4.000 436.240 896.000 436.880 ;
        RECT 4.000 434.840 895.600 436.240 ;
        RECT 4.000 426.040 896.000 434.840 ;
        RECT 4.400 424.640 896.000 426.040 ;
        RECT 4.000 421.960 896.000 424.640 ;
        RECT 4.000 420.560 895.600 421.960 ;
        RECT 4.000 413.800 896.000 420.560 ;
        RECT 4.400 412.400 896.000 413.800 ;
        RECT 4.000 407.680 896.000 412.400 ;
        RECT 4.000 406.280 895.600 407.680 ;
        RECT 4.000 402.240 896.000 406.280 ;
        RECT 4.400 400.840 896.000 402.240 ;
        RECT 4.000 393.400 896.000 400.840 ;
        RECT 4.000 392.000 895.600 393.400 ;
        RECT 4.000 390.000 896.000 392.000 ;
        RECT 4.400 388.600 896.000 390.000 ;
        RECT 4.000 379.120 896.000 388.600 ;
        RECT 4.000 377.760 895.600 379.120 ;
        RECT 4.400 377.720 895.600 377.760 ;
        RECT 4.400 376.360 896.000 377.720 ;
        RECT 4.000 366.200 896.000 376.360 ;
        RECT 4.400 364.840 896.000 366.200 ;
        RECT 4.400 364.800 895.600 364.840 ;
        RECT 4.000 363.440 895.600 364.800 ;
        RECT 4.000 353.960 896.000 363.440 ;
        RECT 4.400 352.560 896.000 353.960 ;
        RECT 4.000 350.560 896.000 352.560 ;
        RECT 4.000 349.160 895.600 350.560 ;
        RECT 4.000 341.720 896.000 349.160 ;
        RECT 4.400 340.320 896.000 341.720 ;
        RECT 4.000 336.280 896.000 340.320 ;
        RECT 4.000 334.880 895.600 336.280 ;
        RECT 4.000 330.160 896.000 334.880 ;
        RECT 4.400 328.760 896.000 330.160 ;
        RECT 4.000 322.000 896.000 328.760 ;
        RECT 4.000 320.600 895.600 322.000 ;
        RECT 4.000 317.920 896.000 320.600 ;
        RECT 4.400 316.520 896.000 317.920 ;
        RECT 4.000 307.720 896.000 316.520 ;
        RECT 4.000 306.360 895.600 307.720 ;
        RECT 4.400 306.320 895.600 306.360 ;
        RECT 4.400 304.960 896.000 306.320 ;
        RECT 4.000 294.120 896.000 304.960 ;
        RECT 4.400 293.440 896.000 294.120 ;
        RECT 4.400 292.720 895.600 293.440 ;
        RECT 4.000 292.040 895.600 292.720 ;
        RECT 4.000 281.880 896.000 292.040 ;
        RECT 4.400 280.480 896.000 281.880 ;
        RECT 4.000 279.160 896.000 280.480 ;
        RECT 4.000 277.760 895.600 279.160 ;
        RECT 4.000 270.320 896.000 277.760 ;
        RECT 4.400 268.920 896.000 270.320 ;
        RECT 4.000 264.880 896.000 268.920 ;
        RECT 4.000 263.480 895.600 264.880 ;
        RECT 4.000 258.080 896.000 263.480 ;
        RECT 4.400 256.680 896.000 258.080 ;
        RECT 4.000 250.600 896.000 256.680 ;
        RECT 4.000 249.200 895.600 250.600 ;
        RECT 4.000 245.840 896.000 249.200 ;
        RECT 4.400 244.440 896.000 245.840 ;
        RECT 4.000 236.320 896.000 244.440 ;
        RECT 4.000 234.920 895.600 236.320 ;
        RECT 4.000 234.280 896.000 234.920 ;
        RECT 4.400 232.880 896.000 234.280 ;
        RECT 4.000 222.040 896.000 232.880 ;
        RECT 4.400 220.640 895.600 222.040 ;
        RECT 4.000 209.800 896.000 220.640 ;
        RECT 4.400 208.400 896.000 209.800 ;
        RECT 4.000 207.760 896.000 208.400 ;
        RECT 4.000 206.360 895.600 207.760 ;
        RECT 4.000 198.240 896.000 206.360 ;
        RECT 4.400 196.840 896.000 198.240 ;
        RECT 4.000 193.480 896.000 196.840 ;
        RECT 4.000 192.080 895.600 193.480 ;
        RECT 4.000 186.000 896.000 192.080 ;
        RECT 4.400 184.600 896.000 186.000 ;
        RECT 4.000 179.200 896.000 184.600 ;
        RECT 4.000 177.800 895.600 179.200 ;
        RECT 4.000 173.760 896.000 177.800 ;
        RECT 4.400 172.360 896.000 173.760 ;
        RECT 4.000 164.920 896.000 172.360 ;
        RECT 4.000 163.520 895.600 164.920 ;
        RECT 4.000 162.200 896.000 163.520 ;
        RECT 4.400 160.800 896.000 162.200 ;
        RECT 4.000 150.640 896.000 160.800 ;
        RECT 4.000 149.960 895.600 150.640 ;
        RECT 4.400 149.240 895.600 149.960 ;
        RECT 4.400 148.560 896.000 149.240 ;
        RECT 4.000 138.400 896.000 148.560 ;
        RECT 4.400 137.000 896.000 138.400 ;
        RECT 4.000 136.360 896.000 137.000 ;
        RECT 4.000 134.960 895.600 136.360 ;
        RECT 4.000 126.160 896.000 134.960 ;
        RECT 4.400 124.760 896.000 126.160 ;
        RECT 4.000 122.080 896.000 124.760 ;
        RECT 4.000 120.680 895.600 122.080 ;
        RECT 4.000 113.920 896.000 120.680 ;
        RECT 4.400 112.520 896.000 113.920 ;
        RECT 4.000 107.800 896.000 112.520 ;
        RECT 4.000 106.400 895.600 107.800 ;
        RECT 4.000 102.360 896.000 106.400 ;
        RECT 4.400 100.960 896.000 102.360 ;
        RECT 4.000 93.520 896.000 100.960 ;
        RECT 4.000 92.120 895.600 93.520 ;
        RECT 4.000 90.120 896.000 92.120 ;
        RECT 4.400 88.720 896.000 90.120 ;
        RECT 4.000 79.240 896.000 88.720 ;
        RECT 4.000 77.880 895.600 79.240 ;
        RECT 4.400 77.840 895.600 77.880 ;
        RECT 4.400 76.480 896.000 77.840 ;
        RECT 4.000 66.320 896.000 76.480 ;
        RECT 4.400 64.960 896.000 66.320 ;
        RECT 4.400 64.920 895.600 64.960 ;
        RECT 4.000 63.560 895.600 64.920 ;
        RECT 4.000 54.080 896.000 63.560 ;
        RECT 4.400 52.680 896.000 54.080 ;
        RECT 4.000 50.680 896.000 52.680 ;
        RECT 4.000 49.280 895.600 50.680 ;
        RECT 4.000 41.840 896.000 49.280 ;
        RECT 4.400 40.440 896.000 41.840 ;
        RECT 4.000 36.400 896.000 40.440 ;
        RECT 4.000 35.000 895.600 36.400 ;
        RECT 4.000 30.280 896.000 35.000 ;
        RECT 4.400 28.880 896.000 30.280 ;
        RECT 4.000 22.120 896.000 28.880 ;
        RECT 4.000 20.720 895.600 22.120 ;
        RECT 4.000 18.040 896.000 20.720 ;
        RECT 4.400 16.640 896.000 18.040 ;
        RECT 4.000 7.840 896.000 16.640 ;
        RECT 4.000 6.480 895.600 7.840 ;
        RECT 4.400 6.440 895.600 6.480 ;
        RECT 4.400 5.630 896.000 6.440 ;
      LAYER met4 ;
        RECT 227.535 10.240 251.040 273.185 ;
        RECT 253.440 10.480 254.340 273.185 ;
        RECT 256.740 10.480 257.640 273.185 ;
        RECT 260.040 10.480 260.940 273.185 ;
        RECT 263.340 10.480 323.545 273.185 ;
        RECT 253.440 10.240 323.545 10.480 ;
        RECT 227.535 6.295 323.545 10.240 ;
  END
END subservient
END LIBRARY

