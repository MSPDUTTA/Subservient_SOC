VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO subservient
  CLASS BLOCK ;
  FOREIGN subservient ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN i_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END i_clk
  PIN i_debug_mode
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 596.000 14.170 600.000 ;
    END
  END i_debug_mode
  PIN i_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END i_rst
  PIN i_sram_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END i_sram_rdata[0]
  PIN i_sram_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 596.000 154.470 600.000 ;
    END
  END i_sram_rdata[1]
  PIN i_sram_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END i_sram_rdata[2]
  PIN i_sram_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END i_sram_rdata[3]
  PIN i_sram_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END i_sram_rdata[4]
  PIN i_sram_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 0.000 322.830 4.000 ;
    END
  END i_sram_rdata[5]
  PIN i_sram_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 241.440 900.000 242.040 ;
    END
  END i_sram_rdata[6]
  PIN i_sram_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 299.240 900.000 299.840 ;
    END
  END i_sram_rdata[7]
  PIN i_wb_dbg_adr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END i_wb_dbg_adr[0]
  PIN i_wb_dbg_adr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.730 0.000 499.010 4.000 ;
    END
  END i_wb_dbg_adr[10]
  PIN i_wb_dbg_adr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.080 4.000 308.680 ;
    END
  END i_wb_dbg_adr[11]
  PIN i_wb_dbg_adr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END i_wb_dbg_adr[12]
  PIN i_wb_dbg_adr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 0.000 538.110 4.000 ;
    END
  END i_wb_dbg_adr[13]
  PIN i_wb_dbg_adr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END i_wb_dbg_adr[14]
  PIN i_wb_dbg_adr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.610 0.000 557.890 4.000 ;
    END
  END i_wb_dbg_adr[15]
  PIN i_wb_dbg_adr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END i_wb_dbg_adr[16]
  PIN i_wb_dbg_adr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.030 0.000 616.310 4.000 ;
    END
  END i_wb_dbg_adr[17]
  PIN i_wb_dbg_adr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 596.000 576.750 600.000 ;
    END
  END i_wb_dbg_adr[18]
  PIN i_wb_dbg_adr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.200 4.000 484.800 ;
    END
  END i_wb_dbg_adr[19]
  PIN i_wb_dbg_adr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END i_wb_dbg_adr[1]
  PIN i_wb_dbg_adr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.130 0.000 655.410 4.000 ;
    END
  END i_wb_dbg_adr[20]
  PIN i_wb_dbg_adr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 596.000 604.810 600.000 ;
    END
  END i_wb_dbg_adr[21]
  PIN i_wb_dbg_adr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END i_wb_dbg_adr[22]
  PIN i_wb_dbg_adr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.790 0.000 734.070 4.000 ;
    END
  END i_wb_dbg_adr[23]
  PIN i_wb_dbg_adr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.110 0.000 753.390 4.000 ;
    END
  END i_wb_dbg_adr[24]
  PIN i_wb_dbg_adr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 512.080 900.000 512.680 ;
    END
  END i_wb_dbg_adr[25]
  PIN i_wb_dbg_adr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 596.000 745.570 600.000 ;
    END
  END i_wb_dbg_adr[26]
  PIN i_wb_dbg_adr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 570.560 900.000 571.160 ;
    END
  END i_wb_dbg_adr[27]
  PIN i_wb_dbg_adr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.470 596.000 829.750 600.000 ;
    END
  END i_wb_dbg_adr[28]
  PIN i_wb_dbg_adr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.990 0.000 812.270 4.000 ;
    END
  END i_wb_dbg_adr[29]
  PIN i_wb_dbg_adr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END i_wb_dbg_adr[2]
  PIN i_wb_dbg_adr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.280 4.000 590.880 ;
    END
  END i_wb_dbg_adr[30]
  PIN i_wb_dbg_adr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.190 0.000 890.470 4.000 ;
    END
  END i_wb_dbg_adr[31]
  PIN i_wb_dbg_adr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 86.400 900.000 87.000 ;
    END
  END i_wb_dbg_adr[3]
  PIN i_wb_dbg_adr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END i_wb_dbg_adr[4]
  PIN i_wb_dbg_adr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END i_wb_dbg_adr[5]
  PIN i_wb_dbg_adr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END i_wb_dbg_adr[6]
  PIN i_wb_dbg_adr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 318.960 900.000 319.560 ;
    END
  END i_wb_dbg_adr[7]
  PIN i_wb_dbg_adr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 357.720 900.000 358.320 ;
    END
  END i_wb_dbg_adr[8]
  PIN i_wb_dbg_adr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.630 0.000 459.910 4.000 ;
    END
  END i_wb_dbg_adr[9]
  PIN i_wb_dbg_dat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 596.000 98.350 600.000 ;
    END
  END i_wb_dbg_dat[0]
  PIN i_wb_dbg_dat[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.720 4.000 273.320 ;
    END
  END i_wb_dbg_dat[10]
  PIN i_wb_dbg_dat[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 4.000 ;
    END
  END i_wb_dbg_dat[11]
  PIN i_wb_dbg_dat[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 396.480 900.000 397.080 ;
    END
  END i_wb_dbg_dat[12]
  PIN i_wb_dbg_dat[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END i_wb_dbg_dat[13]
  PIN i_wb_dbg_dat[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END i_wb_dbg_dat[14]
  PIN i_wb_dbg_dat[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END i_wb_dbg_dat[15]
  PIN i_wb_dbg_dat[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.160 4.000 431.760 ;
    END
  END i_wb_dbg_dat[16]
  PIN i_wb_dbg_dat[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 596.000 548.230 600.000 ;
    END
  END i_wb_dbg_dat[17]
  PIN i_wb_dbg_dat[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END i_wb_dbg_dat[18]
  PIN i_wb_dbg_dat[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 473.320 900.000 473.920 ;
    END
  END i_wb_dbg_dat[19]
  PIN i_wb_dbg_dat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 596.000 182.530 600.000 ;
    END
  END i_wb_dbg_dat[1]
  PIN i_wb_dbg_dat[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.880 4.000 502.480 ;
    END
  END i_wb_dbg_dat[20]
  PIN i_wb_dbg_dat[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.590 596.000 632.870 600.000 ;
    END
  END i_wb_dbg_dat[21]
  PIN i_wb_dbg_dat[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.690 0.000 694.970 4.000 ;
    END
  END i_wb_dbg_dat[22]
  PIN i_wb_dbg_dat[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 493.040 900.000 493.640 ;
    END
  END i_wb_dbg_dat[23]
  PIN i_wb_dbg_dat[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 596.000 660.930 600.000 ;
    END
  END i_wb_dbg_dat[24]
  PIN i_wb_dbg_dat[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 531.800 900.000 532.400 ;
    END
  END i_wb_dbg_dat[25]
  PIN i_wb_dbg_dat[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 0.000 773.170 4.000 ;
    END
  END i_wb_dbg_dat[26]
  PIN i_wb_dbg_dat[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.350 596.000 773.630 600.000 ;
    END
  END i_wb_dbg_dat[27]
  PIN i_wb_dbg_dat[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 0.000 792.490 4.000 ;
    END
  END i_wb_dbg_dat[28]
  PIN i_wb_dbg_dat[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.310 0.000 831.590 4.000 ;
    END
  END i_wb_dbg_dat[29]
  PIN i_wb_dbg_dat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END i_wb_dbg_dat[2]
  PIN i_wb_dbg_dat[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.090 0.000 851.370 4.000 ;
    END
  END i_wb_dbg_dat[30]
  PIN i_wb_dbg_dat[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.590 596.000 885.870 600.000 ;
    END
  END i_wb_dbg_dat[31]
  PIN i_wb_dbg_dat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 106.120 900.000 106.720 ;
    END
  END i_wb_dbg_dat[3]
  PIN i_wb_dbg_dat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 0.000 303.510 4.000 ;
    END
  END i_wb_dbg_dat[4]
  PIN i_wb_dbg_dat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 596.000 323.290 600.000 ;
    END
  END i_wb_dbg_dat[5]
  PIN i_wb_dbg_dat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 260.480 900.000 261.080 ;
    END
  END i_wb_dbg_dat[6]
  PIN i_wb_dbg_dat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 596.000 407.930 600.000 ;
    END
  END i_wb_dbg_dat[7]
  PIN i_wb_dbg_dat[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END i_wb_dbg_dat[8]
  PIN i_wb_dbg_dat[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.830 596.000 492.110 600.000 ;
    END
  END i_wb_dbg_dat[9]
  PIN i_wb_dbg_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 9.560 900.000 10.160 ;
    END
  END i_wb_dbg_sel[0]
  PIN i_wb_dbg_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 596.000 211.050 600.000 ;
    END
  END i_wb_dbg_sel[1]
  PIN i_wb_dbg_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 4.000 96.520 ;
    END
  END i_wb_dbg_sel[2]
  PIN i_wb_dbg_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 0.000 244.630 4.000 ;
    END
  END i_wb_dbg_sel[3]
  PIN i_wb_dbg_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 596.000 42.230 600.000 ;
    END
  END i_wb_dbg_stb
  PIN i_wb_dbg_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END i_wb_dbg_we
  PIN o_gpio
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END o_gpio
  PIN o_sram_raddr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END o_sram_raddr[0]
  PIN o_sram_raddr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 596.000 239.110 600.000 ;
    END
  END o_sram_raddr[1]
  PIN o_sram_raddr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 47.640 900.000 48.240 ;
    END
  END o_sram_raddr[2]
  PIN o_sram_raddr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END o_sram_raddr[3]
  PIN o_sram_raddr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 144.880 900.000 145.480 ;
    END
  END o_sram_raddr[4]
  PIN o_sram_raddr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 4.000 ;
    END
  END o_sram_raddr[5]
  PIN o_sram_raddr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 280.200 900.000 280.800 ;
    END
  END o_sram_raddr[6]
  PIN o_sram_raddr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.710 596.000 435.990 600.000 ;
    END
  END o_sram_raddr[7]
  PIN o_sram_raddr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.770 596.000 464.050 600.000 ;
    END
  END o_sram_raddr[8]
  PIN o_sram_ren
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 596.000 70.290 600.000 ;
    END
  END o_sram_ren
  PIN o_sram_waddr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 596.000 126.410 600.000 ;
    END
  END o_sram_waddr[0]
  PIN o_sram_waddr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 596.000 267.170 600.000 ;
    END
  END o_sram_waddr[1]
  PIN o_sram_waddr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END o_sram_waddr[2]
  PIN o_sram_waddr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 125.160 900.000 125.760 ;
    END
  END o_sram_waddr[3]
  PIN o_sram_waddr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 163.920 900.000 164.520 ;
    END
  END o_sram_waddr[4]
  PIN o_sram_waddr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 0.000 381.710 4.000 ;
    END
  END o_sram_waddr[5]
  PIN o_sram_waddr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.000 4.000 202.600 ;
    END
  END o_sram_waddr[6]
  PIN o_sram_waddr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.360 4.000 237.960 ;
    END
  END o_sram_waddr[7]
  PIN o_sram_waddr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 0.000 420.810 4.000 ;
    END
  END o_sram_waddr[8]
  PIN o_sram_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END o_sram_wdata[0]
  PIN o_sram_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 4.000 61.160 ;
    END
  END o_sram_wdata[1]
  PIN o_sram_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 67.360 900.000 67.960 ;
    END
  END o_sram_wdata[2]
  PIN o_sram_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 4.000 131.880 ;
    END
  END o_sram_wdata[3]
  PIN o_sram_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 183.640 900.000 184.240 ;
    END
  END o_sram_wdata[4]
  PIN o_sram_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 596.000 351.350 600.000 ;
    END
  END o_sram_wdata[5]
  PIN o_sram_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END o_sram_wdata[6]
  PIN o_sram_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.750 0.000 401.030 4.000 ;
    END
  END o_sram_wdata[7]
  PIN o_sram_wen
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END o_sram_wen
  PIN o_wb_dbg_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END o_wb_dbg_ack
  PIN o_wb_dbg_rdt[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 28.600 900.000 29.200 ;
    END
  END o_wb_dbg_rdt[0]
  PIN o_wb_dbg_rdt[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 290.400 4.000 291.000 ;
    END
  END o_wb_dbg_rdt[10]
  PIN o_wb_dbg_rdt[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 376.760 900.000 377.360 ;
    END
  END o_wb_dbg_rdt[11]
  PIN o_wb_dbg_rdt[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 415.520 900.000 416.120 ;
    END
  END o_wb_dbg_rdt[12]
  PIN o_wb_dbg_rdt[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 434.560 900.000 435.160 ;
    END
  END o_wb_dbg_rdt[13]
  PIN o_wb_dbg_rdt[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.890 596.000 520.170 600.000 ;
    END
  END o_wb_dbg_rdt[14]
  PIN o_wb_dbg_rdt[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.930 0.000 577.210 4.000 ;
    END
  END o_wb_dbg_rdt[15]
  PIN o_wb_dbg_rdt[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.710 0.000 596.990 4.000 ;
    END
  END o_wb_dbg_rdt[16]
  PIN o_wb_dbg_rdt[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 454.280 900.000 454.880 ;
    END
  END o_wb_dbg_rdt[17]
  PIN o_wb_dbg_rdt[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.520 4.000 467.120 ;
    END
  END o_wb_dbg_rdt[18]
  PIN o_wb_dbg_rdt[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.810 0.000 636.090 4.000 ;
    END
  END o_wb_dbg_rdt[19]
  PIN o_wb_dbg_rdt[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END o_wb_dbg_rdt[1]
  PIN o_wb_dbg_rdt[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.560 4.000 520.160 ;
    END
  END o_wb_dbg_rdt[20]
  PIN o_wb_dbg_rdt[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 0.000 675.190 4.000 ;
    END
  END o_wb_dbg_rdt[21]
  PIN o_wb_dbg_rdt[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.010 0.000 714.290 4.000 ;
    END
  END o_wb_dbg_rdt[22]
  PIN o_wb_dbg_rdt[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.920 4.000 555.520 ;
    END
  END o_wb_dbg_rdt[23]
  PIN o_wb_dbg_rdt[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.710 596.000 688.990 600.000 ;
    END
  END o_wb_dbg_rdt[24]
  PIN o_wb_dbg_rdt[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.770 596.000 717.050 600.000 ;
    END
  END o_wb_dbg_rdt[25]
  PIN o_wb_dbg_rdt[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 550.840 900.000 551.440 ;
    END
  END o_wb_dbg_rdt[26]
  PIN o_wb_dbg_rdt[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.410 596.000 801.690 600.000 ;
    END
  END o_wb_dbg_rdt[27]
  PIN o_wb_dbg_rdt[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.530 596.000 857.810 600.000 ;
    END
  END o_wb_dbg_rdt[28]
  PIN o_wb_dbg_rdt[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 572.600 4.000 573.200 ;
    END
  END o_wb_dbg_rdt[29]
  PIN o_wb_dbg_rdt[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 596.000 295.230 600.000 ;
    END
  END o_wb_dbg_rdt[2]
  PIN o_wb_dbg_rdt[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.410 0.000 870.690 4.000 ;
    END
  END o_wb_dbg_rdt[30]
  PIN o_wb_dbg_rdt[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 589.600 900.000 590.200 ;
    END
  END o_wb_dbg_rdt[31]
  PIN o_wb_dbg_rdt[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END o_wb_dbg_rdt[3]
  PIN o_wb_dbg_rdt[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 202.680 900.000 203.280 ;
    END
  END o_wb_dbg_rdt[4]
  PIN o_wb_dbg_rdt[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 221.720 900.000 222.320 ;
    END
  END o_wb_dbg_rdt[5]
  PIN o_wb_dbg_rdt[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 596.000 379.870 600.000 ;
    END
  END o_wb_dbg_rdt[6]
  PIN o_wb_dbg_rdt[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 338.000 900.000 338.600 ;
    END
  END o_wb_dbg_rdt[7]
  PIN o_wb_dbg_rdt[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 0.000 440.130 4.000 ;
    END
  END o_wb_dbg_rdt[8]
  PIN o_wb_dbg_rdt[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 0.000 479.690 4.000 ;
    END
  END o_wb_dbg_rdt[9]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 587.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 587.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 486.030 894.240 487.630 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 332.850 894.240 334.450 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 179.670 894.240 181.270 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 894.240 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 587.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 587.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 562.620 894.240 564.220 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 409.440 894.240 411.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 256.260 894.240 257.860 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 894.240 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 215.425 11.305 505.855 270.895 ;
      LAYER met1 ;
        RECT 5.520 10.640 894.240 587.760 ;
      LAYER met2 ;
        RECT 9.760 595.720 13.610 596.000 ;
        RECT 14.450 595.720 41.670 596.000 ;
        RECT 42.510 595.720 69.730 596.000 ;
        RECT 70.570 595.720 97.790 596.000 ;
        RECT 98.630 595.720 125.850 596.000 ;
        RECT 126.690 595.720 153.910 596.000 ;
        RECT 154.750 595.720 181.970 596.000 ;
        RECT 182.810 595.720 210.490 596.000 ;
        RECT 211.330 595.720 238.550 596.000 ;
        RECT 239.390 595.720 266.610 596.000 ;
        RECT 267.450 595.720 294.670 596.000 ;
        RECT 295.510 595.720 322.730 596.000 ;
        RECT 323.570 595.720 350.790 596.000 ;
        RECT 351.630 595.720 379.310 596.000 ;
        RECT 380.150 595.720 407.370 596.000 ;
        RECT 408.210 595.720 435.430 596.000 ;
        RECT 436.270 595.720 463.490 596.000 ;
        RECT 464.330 595.720 491.550 596.000 ;
        RECT 492.390 595.720 519.610 596.000 ;
        RECT 520.450 595.720 547.670 596.000 ;
        RECT 548.510 595.720 576.190 596.000 ;
        RECT 577.030 595.720 604.250 596.000 ;
        RECT 605.090 595.720 632.310 596.000 ;
        RECT 633.150 595.720 660.370 596.000 ;
        RECT 661.210 595.720 688.430 596.000 ;
        RECT 689.270 595.720 716.490 596.000 ;
        RECT 717.330 595.720 745.010 596.000 ;
        RECT 745.850 595.720 773.070 596.000 ;
        RECT 773.910 595.720 801.130 596.000 ;
        RECT 801.970 595.720 829.190 596.000 ;
        RECT 830.030 595.720 857.250 596.000 ;
        RECT 858.090 595.720 885.310 596.000 ;
        RECT 886.150 595.720 890.460 596.000 ;
        RECT 9.760 4.280 890.460 595.720 ;
        RECT 10.310 4.000 28.790 4.280 ;
        RECT 29.630 4.000 48.570 4.280 ;
        RECT 49.410 4.000 67.890 4.280 ;
        RECT 68.730 4.000 87.670 4.280 ;
        RECT 88.510 4.000 106.990 4.280 ;
        RECT 107.830 4.000 126.770 4.280 ;
        RECT 127.610 4.000 146.090 4.280 ;
        RECT 146.930 4.000 165.870 4.280 ;
        RECT 166.710 4.000 185.190 4.280 ;
        RECT 186.030 4.000 204.970 4.280 ;
        RECT 205.810 4.000 224.290 4.280 ;
        RECT 225.130 4.000 244.070 4.280 ;
        RECT 244.910 4.000 263.850 4.280 ;
        RECT 264.690 4.000 283.170 4.280 ;
        RECT 284.010 4.000 302.950 4.280 ;
        RECT 303.790 4.000 322.270 4.280 ;
        RECT 323.110 4.000 342.050 4.280 ;
        RECT 342.890 4.000 361.370 4.280 ;
        RECT 362.210 4.000 381.150 4.280 ;
        RECT 381.990 4.000 400.470 4.280 ;
        RECT 401.310 4.000 420.250 4.280 ;
        RECT 421.090 4.000 439.570 4.280 ;
        RECT 440.410 4.000 459.350 4.280 ;
        RECT 460.190 4.000 479.130 4.280 ;
        RECT 479.970 4.000 498.450 4.280 ;
        RECT 499.290 4.000 518.230 4.280 ;
        RECT 519.070 4.000 537.550 4.280 ;
        RECT 538.390 4.000 557.330 4.280 ;
        RECT 558.170 4.000 576.650 4.280 ;
        RECT 577.490 4.000 596.430 4.280 ;
        RECT 597.270 4.000 615.750 4.280 ;
        RECT 616.590 4.000 635.530 4.280 ;
        RECT 636.370 4.000 654.850 4.280 ;
        RECT 655.690 4.000 674.630 4.280 ;
        RECT 675.470 4.000 694.410 4.280 ;
        RECT 695.250 4.000 713.730 4.280 ;
        RECT 714.570 4.000 733.510 4.280 ;
        RECT 734.350 4.000 752.830 4.280 ;
        RECT 753.670 4.000 772.610 4.280 ;
        RECT 773.450 4.000 791.930 4.280 ;
        RECT 792.770 4.000 811.710 4.280 ;
        RECT 812.550 4.000 831.030 4.280 ;
        RECT 831.870 4.000 850.810 4.280 ;
        RECT 851.650 4.000 870.130 4.280 ;
        RECT 870.970 4.000 889.910 4.280 ;
      LAYER met3 ;
        RECT 4.400 590.600 896.000 590.745 ;
        RECT 4.400 589.880 895.600 590.600 ;
        RECT 4.000 589.200 895.600 589.880 ;
        RECT 4.000 573.600 896.000 589.200 ;
        RECT 4.400 572.200 896.000 573.600 ;
        RECT 4.000 571.560 896.000 572.200 ;
        RECT 4.000 570.160 895.600 571.560 ;
        RECT 4.000 555.920 896.000 570.160 ;
        RECT 4.400 554.520 896.000 555.920 ;
        RECT 4.000 551.840 896.000 554.520 ;
        RECT 4.000 550.440 895.600 551.840 ;
        RECT 4.000 538.240 896.000 550.440 ;
        RECT 4.400 536.840 896.000 538.240 ;
        RECT 4.000 532.800 896.000 536.840 ;
        RECT 4.000 531.400 895.600 532.800 ;
        RECT 4.000 520.560 896.000 531.400 ;
        RECT 4.400 519.160 896.000 520.560 ;
        RECT 4.000 513.080 896.000 519.160 ;
        RECT 4.000 511.680 895.600 513.080 ;
        RECT 4.000 502.880 896.000 511.680 ;
        RECT 4.400 501.480 896.000 502.880 ;
        RECT 4.000 494.040 896.000 501.480 ;
        RECT 4.000 492.640 895.600 494.040 ;
        RECT 4.000 485.200 896.000 492.640 ;
        RECT 4.400 483.800 896.000 485.200 ;
        RECT 4.000 474.320 896.000 483.800 ;
        RECT 4.000 472.920 895.600 474.320 ;
        RECT 4.000 467.520 896.000 472.920 ;
        RECT 4.400 466.120 896.000 467.520 ;
        RECT 4.000 455.280 896.000 466.120 ;
        RECT 4.000 453.880 895.600 455.280 ;
        RECT 4.000 449.840 896.000 453.880 ;
        RECT 4.400 448.440 896.000 449.840 ;
        RECT 4.000 435.560 896.000 448.440 ;
        RECT 4.000 434.160 895.600 435.560 ;
        RECT 4.000 432.160 896.000 434.160 ;
        RECT 4.400 430.760 896.000 432.160 ;
        RECT 4.000 416.520 896.000 430.760 ;
        RECT 4.000 415.120 895.600 416.520 ;
        RECT 4.000 414.480 896.000 415.120 ;
        RECT 4.400 413.080 896.000 414.480 ;
        RECT 4.000 397.480 896.000 413.080 ;
        RECT 4.000 396.800 895.600 397.480 ;
        RECT 4.400 396.080 895.600 396.800 ;
        RECT 4.400 395.400 896.000 396.080 ;
        RECT 4.000 379.120 896.000 395.400 ;
        RECT 4.400 377.760 896.000 379.120 ;
        RECT 4.400 377.720 895.600 377.760 ;
        RECT 4.000 376.360 895.600 377.720 ;
        RECT 4.000 361.440 896.000 376.360 ;
        RECT 4.400 360.040 896.000 361.440 ;
        RECT 4.000 358.720 896.000 360.040 ;
        RECT 4.000 357.320 895.600 358.720 ;
        RECT 4.000 343.760 896.000 357.320 ;
        RECT 4.400 342.360 896.000 343.760 ;
        RECT 4.000 339.000 896.000 342.360 ;
        RECT 4.000 337.600 895.600 339.000 ;
        RECT 4.000 326.080 896.000 337.600 ;
        RECT 4.400 324.680 896.000 326.080 ;
        RECT 4.000 319.960 896.000 324.680 ;
        RECT 4.000 318.560 895.600 319.960 ;
        RECT 4.000 309.080 896.000 318.560 ;
        RECT 4.400 307.680 896.000 309.080 ;
        RECT 4.000 300.240 896.000 307.680 ;
        RECT 4.000 298.840 895.600 300.240 ;
        RECT 4.000 291.400 896.000 298.840 ;
        RECT 4.400 290.000 896.000 291.400 ;
        RECT 4.000 281.200 896.000 290.000 ;
        RECT 4.000 279.800 895.600 281.200 ;
        RECT 4.000 273.720 896.000 279.800 ;
        RECT 4.400 272.320 896.000 273.720 ;
        RECT 4.000 261.480 896.000 272.320 ;
        RECT 4.000 260.080 895.600 261.480 ;
        RECT 4.000 256.040 896.000 260.080 ;
        RECT 4.400 254.640 896.000 256.040 ;
        RECT 4.000 242.440 896.000 254.640 ;
        RECT 4.000 241.040 895.600 242.440 ;
        RECT 4.000 238.360 896.000 241.040 ;
        RECT 4.400 236.960 896.000 238.360 ;
        RECT 4.000 222.720 896.000 236.960 ;
        RECT 4.000 221.320 895.600 222.720 ;
        RECT 4.000 220.680 896.000 221.320 ;
        RECT 4.400 219.280 896.000 220.680 ;
        RECT 4.000 203.680 896.000 219.280 ;
        RECT 4.000 203.000 895.600 203.680 ;
        RECT 4.400 202.280 895.600 203.000 ;
        RECT 4.400 201.600 896.000 202.280 ;
        RECT 4.000 185.320 896.000 201.600 ;
        RECT 4.400 184.640 896.000 185.320 ;
        RECT 4.400 183.920 895.600 184.640 ;
        RECT 4.000 183.240 895.600 183.920 ;
        RECT 4.000 167.640 896.000 183.240 ;
        RECT 4.400 166.240 896.000 167.640 ;
        RECT 4.000 164.920 896.000 166.240 ;
        RECT 4.000 163.520 895.600 164.920 ;
        RECT 4.000 149.960 896.000 163.520 ;
        RECT 4.400 148.560 896.000 149.960 ;
        RECT 4.000 145.880 896.000 148.560 ;
        RECT 4.000 144.480 895.600 145.880 ;
        RECT 4.000 132.280 896.000 144.480 ;
        RECT 4.400 130.880 896.000 132.280 ;
        RECT 4.000 126.160 896.000 130.880 ;
        RECT 4.000 124.760 895.600 126.160 ;
        RECT 4.000 114.600 896.000 124.760 ;
        RECT 4.400 113.200 896.000 114.600 ;
        RECT 4.000 107.120 896.000 113.200 ;
        RECT 4.000 105.720 895.600 107.120 ;
        RECT 4.000 96.920 896.000 105.720 ;
        RECT 4.400 95.520 896.000 96.920 ;
        RECT 4.000 87.400 896.000 95.520 ;
        RECT 4.000 86.000 895.600 87.400 ;
        RECT 4.000 79.240 896.000 86.000 ;
        RECT 4.400 77.840 896.000 79.240 ;
        RECT 4.000 68.360 896.000 77.840 ;
        RECT 4.000 66.960 895.600 68.360 ;
        RECT 4.000 61.560 896.000 66.960 ;
        RECT 4.400 60.160 896.000 61.560 ;
        RECT 4.000 48.640 896.000 60.160 ;
        RECT 4.000 47.240 895.600 48.640 ;
        RECT 4.000 43.880 896.000 47.240 ;
        RECT 4.400 42.480 896.000 43.880 ;
        RECT 4.000 29.600 896.000 42.480 ;
        RECT 4.000 28.200 895.600 29.600 ;
        RECT 4.000 26.200 896.000 28.200 ;
        RECT 4.400 24.800 896.000 26.200 ;
        RECT 4.000 10.560 896.000 24.800 ;
        RECT 4.000 9.200 895.600 10.560 ;
        RECT 4.400 9.160 895.600 9.200 ;
        RECT 4.400 8.335 896.000 9.160 ;
      LAYER met4 ;
        RECT 336.095 25.335 336.425 248.705 ;
  END
END subservient
END LIBRARY

